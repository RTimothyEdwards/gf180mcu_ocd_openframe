magic
tech gf180mcuD
magscale 1 10
timestamp 1765161918
<< metal1 >>
rect -244 734 338 854
rect -244 -50 338 70
<< via1 >>
rect 12285 489 12337 657
rect -142 254 -90 422
rect 33 328 85 435
rect 189 281 241 449
rect 491 324 543 467
rect 1612 425 1817 477
rect 1123 225 1175 393
rect 2749 298 2801 466
rect 2877 434 3061 486
rect 3623 429 3828 481
rect 4765 289 4817 457
rect 4893 434 5077 486
rect 5297 328 5349 435
rect 5453 278 5505 446
rect 5880 423 6064 475
rect 7005 292 7057 460
rect 7133 434 7317 486
rect 7666 424 7850 476
rect 8797 295 8849 463
rect 8925 435 9109 487
rect 9686 426 9870 478
rect 10813 290 10865 458
rect 10940 434 11124 486
rect 11427 347 11588 399
rect 11718 347 11879 399
rect 11952 278 12004 446
rect 12626 327 12678 495
<< metal2 >>
rect 2747 654 2803 670
rect 1119 542 1179 560
rect 488 467 546 487
rect -145 422 -86 441
rect -145 254 -142 422
rect -90 254 -86 422
rect -145 206 -86 254
rect 31 435 87 450
rect 31 328 33 435
rect 85 328 87 435
rect 31 206 87 328
rect 185 449 244 464
rect 185 318 189 449
rect 241 318 244 449
rect 488 430 491 467
rect 543 430 546 467
rect 488 324 491 374
rect 543 324 546 374
rect 488 308 546 324
rect 1119 393 1179 486
rect 1594 477 1835 480
rect 1594 425 1612 477
rect 1817 425 1835 477
rect 1594 423 1835 425
rect 2747 466 2803 598
rect 4763 654 4819 667
rect 2958 542 3018 559
rect 185 225 244 262
rect 1119 225 1123 393
rect 1175 225 1179 393
rect 1119 208 1179 225
rect -162 150 -145 206
rect -86 150 -67 206
rect 31 121 87 150
rect 1637 206 1693 423
rect 2747 298 2749 466
rect 2801 298 2803 466
rect 2861 486 2958 490
rect 3018 486 3077 490
rect 2861 434 2877 486
rect 3061 434 3077 486
rect 2861 431 3077 434
rect 3603 481 3847 484
rect 2958 430 3018 431
rect 3603 429 3623 481
rect 3828 429 3847 481
rect 3603 426 3847 429
rect 4763 457 4819 598
rect 5293 654 5353 667
rect 2747 285 2803 298
rect 3659 318 3715 426
rect 4763 289 4765 457
rect 4817 289 4819 457
rect 4881 486 5090 489
rect 4881 434 4893 486
rect 5077 434 5090 486
rect 4881 432 5090 434
rect 5293 435 5353 598
rect 10970 654 11026 666
rect 4980 430 5037 432
rect 4980 357 5037 374
rect 5293 328 5297 435
rect 5349 328 5353 435
rect 5293 304 5353 328
rect 5450 542 5508 565
rect 7191 542 7247 564
rect 5450 446 5508 486
rect 7119 486 7191 489
rect 7681 542 7737 557
rect 7247 486 7331 489
rect 4763 275 4819 289
rect 5450 278 5453 446
rect 5505 278 5508 446
rect 5863 475 6081 478
rect 5863 423 5880 475
rect 6064 423 6081 475
rect 5863 420 6081 423
rect 7002 460 7060 473
rect 7002 430 7005 460
rect 7057 430 7060 460
rect 7119 434 7133 486
rect 7317 434 7331 486
rect 7681 479 7737 486
rect 8913 487 9123 490
rect 10970 489 11026 598
rect 12282 657 12340 669
rect 12282 654 12285 657
rect 12337 654 12340 657
rect 11949 542 12006 553
rect 7119 432 7331 434
rect 7653 476 7865 479
rect 5450 262 5508 278
rect 3659 250 3715 262
rect 1637 136 1693 150
rect 5882 94 5938 420
rect 7653 424 7666 476
rect 7850 424 7865 476
rect 7653 422 7865 424
rect 8795 463 8851 477
rect 8795 430 8797 463
rect 8849 430 8851 463
rect 8913 435 8925 487
rect 9109 435 9123 487
rect 10928 486 11137 489
rect 8913 432 9123 435
rect 9664 478 9889 481
rect 7002 292 7005 374
rect 7057 292 7060 374
rect 7002 274 7060 292
rect 8795 295 8797 374
rect 8849 295 8851 374
rect 8795 246 8851 295
rect 9011 318 9067 432
rect 9664 426 9686 478
rect 9870 426 9889 478
rect 9664 423 9889 426
rect 10810 458 10868 472
rect 10810 430 10813 458
rect 10865 430 10868 458
rect 10928 434 10940 486
rect 11124 434 11137 486
rect 10928 431 11137 434
rect 11949 446 12006 486
rect 12282 489 12285 598
rect 12337 489 12340 598
rect 12282 477 12340 489
rect 12624 495 12680 516
rect 9011 240 9067 262
rect 9694 318 9750 423
rect 10810 290 10813 374
rect 10865 290 10868 374
rect 11411 399 11605 403
rect 11411 347 11427 399
rect 11588 347 11605 399
rect 11411 344 11605 347
rect 11706 399 11892 401
rect 11706 347 11718 399
rect 11879 347 11892 399
rect 11706 345 11892 347
rect 10810 276 10868 290
rect 11433 318 11489 344
rect 9694 251 9750 262
rect 11433 251 11489 262
rect 11770 94 11826 345
rect 11949 278 11952 446
rect 12004 278 12006 446
rect 11949 262 12006 278
rect 12624 327 12626 495
rect 12678 327 12680 495
rect 12624 94 12680 327
rect 5869 38 5882 94
rect 5938 38 5954 94
rect 11757 38 11770 94
rect 11826 38 11839 94
rect 12624 23 12680 38
<< via2 >>
rect 2747 598 2803 654
rect 185 281 189 318
rect 189 281 241 318
rect 241 281 244 318
rect 488 374 491 430
rect 491 374 543 430
rect 543 374 546 430
rect 1119 486 1179 542
rect 4763 598 4819 654
rect 185 262 244 281
rect -145 150 -86 206
rect 31 150 87 206
rect 2958 486 3018 542
rect 5293 598 5353 654
rect 3659 262 3715 318
rect 10970 598 11026 654
rect 4980 374 5037 430
rect 5450 486 5508 542
rect 7191 486 7247 542
rect 7681 486 7737 542
rect 12282 598 12285 654
rect 12285 598 12337 654
rect 12337 598 12340 654
rect 1637 150 1693 206
rect 7002 374 7005 430
rect 7005 374 7057 430
rect 7057 374 7060 430
rect 8795 374 8797 430
rect 8797 374 8849 430
rect 8849 374 8851 430
rect 11949 486 12006 542
rect 9011 262 9067 318
rect 9694 262 9750 318
rect 10810 374 10813 430
rect 10813 374 10865 430
rect 10865 374 10868 430
rect 11433 262 11489 318
rect 5882 38 5938 94
rect 11770 38 11826 94
rect 12624 38 12680 94
<< metal3 >>
rect 2718 598 2747 654
rect 2803 598 4763 654
rect 4819 598 5293 654
rect 5353 598 5391 654
rect 10948 598 10970 654
rect 11026 598 12282 654
rect 12340 598 12362 654
rect 1091 486 1119 542
rect 1179 486 2958 542
rect 3018 486 3043 542
rect 5418 486 5450 542
rect 5508 486 7191 542
rect 7247 486 7348 542
rect 7667 486 7681 542
rect 7737 486 11949 542
rect 12006 486 12032 542
rect 456 374 488 430
rect 546 374 4980 430
rect 5037 374 5251 430
rect 5656 374 7002 430
rect 7060 374 8795 430
rect 8851 374 10810 430
rect 10868 374 10901 430
rect 5195 318 5251 374
rect 160 262 185 318
rect 244 262 3659 318
rect 3715 262 3743 318
rect 5195 262 9011 318
rect 9067 262 9093 318
rect 9677 262 9694 318
rect 9750 262 11433 318
rect 11489 262 12953 318
rect -442 150 -145 206
rect -86 150 31 206
rect 87 150 1637 206
rect 1693 150 12951 206
rect -442 38 5882 94
rect 5938 38 11770 94
rect 11826 38 12624 94
rect 12680 38 12949 94
use gf180mcu_as_sc_mcu7t3v3__tieh_4  const1 $PDKPATH/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532550
transform 1 0 12076 0 1 10
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  ctrlen0 $PDKPATH/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751740063
transform 1 0 11292 0 1 10
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_4  delaybuf0 $PDKPATH/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751558652
transform 1 0 428 0 1 10
box -86 -86 1094 870
use gf180mcu_as_sc_mcu7t3v3__invz_2  delayen0 $PDKPATH/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1764933398
transform 1 0 5692 0 1 10
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__invz_2  delayen1
timestamp 1764933398
transform 1 0 1436 0 1 10
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__invz_2  delayenb0
timestamp 1764933398
transform 1 0 7484 0 1 10
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__invz_2  delayenb1
timestamp 1764933398
transform 1 0 3452 0 1 10
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  delayint0 $PDKPATH/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532043
transform 1 0 5244 0 1 10
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  gf180mcu_as_sc_mcu7t3v3__diode_2_0 $PDKPATH/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532392
transform -1 0 12748 0 1 10
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  gf180mcu_as_sc_mcu7t3v3__diode_2_1
timestamp 1751532392
transform -1 0 -20 0 1 10
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  gf180mcu_as_sc_mcu7t3v3__tap_2_0 $PDKPATH/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1759751540
transform -1 0 -244 0 1 10
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  gf180mcu_as_sc_mcu7t3v3__tap_2_1
timestamp 1759751540
transform -1 0 12972 0 1 10
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  gf180mcu_as_sc_mcu7t3v3__tap_2_2
timestamp 1759751540
transform 1 0 3228 0 1 10
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  gf180mcu_as_sc_mcu7t3v3__tap_2_3
timestamp 1759751540
transform 1 0 9276 0 1 10
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__invz_2  reseten0
timestamp 1764933398
transform 1 0 9500 0 1 10
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  trim1bar
timestamp 1751532043
transform 1 0 -20 0 1 10
box -86 -86 534 870
<< labels >>
flabel metal3 724 374 782 430 0 FreeSans 448 0 0 0 in
port 3 nsew
flabel metal3 1274 262 1334 318 0 FreeSans 448 0 0 0 trim1b
flabel metal3 3206 598 3267 654 0 FreeSans 448 0 0 0 d1
flabel metal3 1268 486 1328 542 0 FreeSans 448 0 0 0 d0
flabel metal3 5527 486 5581 542 0 FreeSans 448 0 0 0 d2
flabel metal3 6733 374 6791 430 0 FreeSans 448 0 0 0 out
port 7 nsew
flabel metal3 11667 486 11725 542 0 FreeSans 448 0 0 0 ctrl0b
flabel metal3 11812 598 11869 654 0 FreeSans 448 0 0 0 one
flabel metal1 -244 734 338 854 0 FreeSans 480 0 0 0 vdd
port 1 nsew
flabel metal1 -244 -50 338 70 0 FreeSans 480 0 0 0 vss
port 2 nsew
flabel metal3 12891 262 12953 318 0 FreeSans 448 0 0 0 reset
port 6 nsew
flabel metal3 -442 38 -387 94 0 FreeSans 448 0 0 0 trim[0]
port 4 nsew
flabel metal3 -442 150 -387 206 0 FreeSans 448 0 0 0 trim[1]
port 5 nsew
<< end >>
