magic
tech gf180mcuD
magscale 1 10
timestamp 1764170769
<< metal1 >>
rect 12323 133 14910 185
rect 15076 133 15452 185
rect 12323 35 15270 87
rect 15436 35 15452 87
<< via1 >>
rect 14910 133 15076 185
rect 15270 35 15436 87
<< metal2 >>
rect 12368 0 12444 232
rect 13241 0 13317 232
rect 15089 187 15145 232
rect 14898 185 15145 187
rect 14898 133 14910 185
rect 15076 133 15145 185
rect 14898 131 15145 133
rect 15089 0 15145 131
rect 15201 89 15257 232
rect 15201 87 15448 89
rect 15201 35 15270 87
rect 15436 35 15448 87
rect 15201 33 15448 35
rect 15201 0 15257 33
<< end >>
