magic
tech gf180mcuD
magscale 1 10
timestamp 1765936290
<< psubdiff >>
rect 0 69943 2000 69968
rect 0 69888 179 69943
rect 0 13160 25 69888
rect 71 69803 179 69888
rect 1823 69888 2000 69943
rect 1823 69803 1929 69888
rect 71 69778 1929 69803
rect 71 13287 93 69778
rect 1907 13287 1929 69778
rect 71 13262 1929 13287
rect 71 13160 179 13262
rect 0 13122 179 13160
rect 1823 13160 1929 13262
rect 1975 13160 2000 69888
rect 1823 13122 2000 13160
rect 0 13097 2000 13122
<< psubdiffcont >>
rect 25 13160 71 69888
rect 179 69803 1823 69943
rect 179 13122 1823 13262
rect 1929 13160 1975 69888
<< metal1 >>
rect -32 69943 2032 69957
rect -32 69888 179 69943
rect -32 13160 25 69888
rect 71 69803 179 69888
rect 1823 69888 2032 69943
rect 1823 69803 1929 69888
rect 71 69789 1929 69803
rect 71 64896 82 69789
rect 1918 64896 1929 69789
rect 71 64884 282 64896
rect 71 64832 94 64884
rect 146 64832 218 64884
rect 270 64832 282 64884
rect 71 64760 282 64832
rect 71 64708 94 64760
rect 146 64708 218 64760
rect 270 64708 282 64760
rect 71 64636 282 64708
rect 71 64584 94 64636
rect 146 64584 218 64636
rect 270 64584 282 64636
rect 71 64512 282 64584
rect 71 64460 94 64512
rect 146 64460 218 64512
rect 270 64460 282 64512
rect 71 64388 282 64460
rect 71 64336 94 64388
rect 146 64336 218 64388
rect 270 64336 282 64388
rect 71 64264 282 64336
rect 71 64212 94 64264
rect 146 64212 218 64264
rect 270 64212 282 64264
rect 71 64140 282 64212
rect 71 64088 94 64140
rect 146 64088 218 64140
rect 270 64088 282 64140
rect 71 64016 282 64088
rect 71 63964 94 64016
rect 146 63964 218 64016
rect 270 63964 282 64016
rect 71 63892 282 63964
rect 71 63840 94 63892
rect 146 63840 218 63892
rect 270 63840 282 63892
rect 71 63768 282 63840
rect 71 63716 94 63768
rect 146 63716 218 63768
rect 270 63716 282 63768
rect 71 63704 282 63716
rect 1718 64884 1929 64896
rect 1718 64832 1730 64884
rect 1782 64832 1854 64884
rect 1906 64832 1929 64884
rect 1718 64760 1929 64832
rect 1718 64708 1730 64760
rect 1782 64708 1854 64760
rect 1906 64708 1929 64760
rect 1718 64636 1929 64708
rect 1718 64584 1730 64636
rect 1782 64584 1854 64636
rect 1906 64584 1929 64636
rect 1718 64512 1929 64584
rect 1718 64460 1730 64512
rect 1782 64460 1854 64512
rect 1906 64460 1929 64512
rect 1718 64388 1929 64460
rect 1718 64336 1730 64388
rect 1782 64336 1854 64388
rect 1906 64336 1929 64388
rect 1718 64264 1929 64336
rect 1718 64212 1730 64264
rect 1782 64212 1854 64264
rect 1906 64212 1929 64264
rect 1718 64140 1929 64212
rect 1718 64088 1730 64140
rect 1782 64088 1854 64140
rect 1906 64088 1929 64140
rect 1718 64016 1929 64088
rect 1718 63964 1730 64016
rect 1782 63964 1854 64016
rect 1906 63964 1929 64016
rect 1718 63892 1929 63964
rect 1718 63840 1730 63892
rect 1782 63840 1854 63892
rect 1906 63840 1929 63892
rect 1718 63768 1929 63840
rect 1718 63716 1730 63768
rect 1782 63716 1854 63768
rect 1906 63716 1929 63768
rect 1718 63704 1929 63716
rect 71 50497 82 63704
rect 1918 50497 1929 63704
rect 71 50485 282 50497
rect 71 50433 94 50485
rect 146 50433 218 50485
rect 270 50433 282 50485
rect 71 50361 282 50433
rect 71 50309 94 50361
rect 146 50309 218 50361
rect 270 50309 282 50361
rect 71 50237 282 50309
rect 71 50185 94 50237
rect 146 50185 218 50237
rect 270 50185 282 50237
rect 71 50113 282 50185
rect 71 50061 94 50113
rect 146 50061 218 50113
rect 270 50061 282 50113
rect 71 49989 282 50061
rect 71 49937 94 49989
rect 146 49937 218 49989
rect 270 49937 282 49989
rect 71 49865 282 49937
rect 71 49813 94 49865
rect 146 49813 218 49865
rect 270 49813 282 49865
rect 71 49741 282 49813
rect 71 49689 94 49741
rect 146 49689 218 49741
rect 270 49689 282 49741
rect 71 49617 282 49689
rect 71 49565 94 49617
rect 146 49565 218 49617
rect 270 49565 282 49617
rect 71 49493 282 49565
rect 71 49441 94 49493
rect 146 49441 218 49493
rect 270 49441 282 49493
rect 71 49369 282 49441
rect 71 49317 94 49369
rect 146 49317 218 49369
rect 270 49317 282 49369
rect 71 49305 282 49317
rect 1718 50485 1929 50497
rect 1718 50433 1730 50485
rect 1782 50433 1854 50485
rect 1906 50433 1929 50485
rect 1718 50361 1929 50433
rect 1718 50309 1730 50361
rect 1782 50309 1854 50361
rect 1906 50309 1929 50361
rect 1718 50237 1929 50309
rect 1718 50185 1730 50237
rect 1782 50185 1854 50237
rect 1906 50185 1929 50237
rect 1718 50113 1929 50185
rect 1718 50061 1730 50113
rect 1782 50061 1854 50113
rect 1906 50061 1929 50113
rect 1718 49989 1929 50061
rect 1718 49937 1730 49989
rect 1782 49937 1854 49989
rect 1906 49937 1929 49989
rect 1718 49865 1929 49937
rect 1718 49813 1730 49865
rect 1782 49813 1854 49865
rect 1906 49813 1929 49865
rect 1718 49741 1929 49813
rect 1718 49689 1730 49741
rect 1782 49689 1854 49741
rect 1906 49689 1929 49741
rect 1718 49617 1929 49689
rect 1718 49565 1730 49617
rect 1782 49565 1854 49617
rect 1906 49565 1929 49617
rect 1718 49493 1929 49565
rect 1718 49441 1730 49493
rect 1782 49441 1854 49493
rect 1906 49441 1929 49493
rect 1718 49369 1929 49441
rect 1718 49317 1730 49369
rect 1782 49317 1854 49369
rect 1906 49317 1929 49369
rect 1718 49305 1929 49317
rect 71 13276 82 49305
rect 1918 13276 1929 49305
rect 71 13262 1929 13276
rect 71 13160 179 13262
rect -32 13122 179 13160
rect 1823 13160 1929 13262
rect 1975 13160 2032 69888
rect 1823 13122 2032 13160
rect -32 13108 2032 13122
<< via1 >>
rect 94 64832 146 64884
rect 218 64832 270 64884
rect 94 64708 146 64760
rect 218 64708 270 64760
rect 94 64584 146 64636
rect 218 64584 270 64636
rect 94 64460 146 64512
rect 218 64460 270 64512
rect 94 64336 146 64388
rect 218 64336 270 64388
rect 94 64212 146 64264
rect 218 64212 270 64264
rect 94 64088 146 64140
rect 218 64088 270 64140
rect 94 63964 146 64016
rect 218 63964 270 64016
rect 94 63840 146 63892
rect 218 63840 270 63892
rect 94 63716 146 63768
rect 218 63716 270 63768
rect 1730 64832 1782 64884
rect 1854 64832 1906 64884
rect 1730 64708 1782 64760
rect 1854 64708 1906 64760
rect 1730 64584 1782 64636
rect 1854 64584 1906 64636
rect 1730 64460 1782 64512
rect 1854 64460 1906 64512
rect 1730 64336 1782 64388
rect 1854 64336 1906 64388
rect 1730 64212 1782 64264
rect 1854 64212 1906 64264
rect 1730 64088 1782 64140
rect 1854 64088 1906 64140
rect 1730 63964 1782 64016
rect 1854 63964 1906 64016
rect 1730 63840 1782 63892
rect 1854 63840 1906 63892
rect 1730 63716 1782 63768
rect 1854 63716 1906 63768
rect 94 50433 146 50485
rect 218 50433 270 50485
rect 94 50309 146 50361
rect 218 50309 270 50361
rect 94 50185 146 50237
rect 218 50185 270 50237
rect 94 50061 146 50113
rect 218 50061 270 50113
rect 94 49937 146 49989
rect 218 49937 270 49989
rect 94 49813 146 49865
rect 218 49813 270 49865
rect 94 49689 146 49741
rect 218 49689 270 49741
rect 94 49565 146 49617
rect 218 49565 270 49617
rect 94 49441 146 49493
rect 218 49441 270 49493
rect 94 49317 146 49369
rect 218 49317 270 49369
rect 1730 50433 1782 50485
rect 1854 50433 1906 50485
rect 1730 50309 1782 50361
rect 1854 50309 1906 50361
rect 1730 50185 1782 50237
rect 1854 50185 1906 50237
rect 1730 50061 1782 50113
rect 1854 50061 1906 50113
rect 1730 49937 1782 49989
rect 1854 49937 1906 49989
rect 1730 49813 1782 49865
rect 1854 49813 1906 49865
rect 1730 49689 1782 49741
rect 1854 49689 1906 49741
rect 1730 49565 1782 49617
rect 1854 49565 1906 49617
rect 1730 49441 1782 49493
rect 1854 49441 1906 49493
rect 1730 49317 1782 49369
rect 1854 49317 1906 49369
<< metal2 >>
rect 0 64886 282 69054
rect 0 64830 92 64886
rect 148 64830 216 64886
rect 272 64830 282 64886
rect 0 64762 282 64830
rect 0 64706 92 64762
rect 148 64706 216 64762
rect 272 64706 282 64762
rect 0 64638 282 64706
rect 0 64582 92 64638
rect 148 64582 216 64638
rect 272 64582 282 64638
rect 0 64514 282 64582
rect 0 64458 92 64514
rect 148 64458 216 64514
rect 272 64458 282 64514
rect 0 64390 282 64458
rect 0 64334 92 64390
rect 148 64334 216 64390
rect 272 64334 282 64390
rect 0 64266 282 64334
rect 0 64210 92 64266
rect 148 64210 216 64266
rect 272 64210 282 64266
rect 0 64142 282 64210
rect 0 64086 92 64142
rect 148 64086 216 64142
rect 272 64086 282 64142
rect 0 64018 282 64086
rect 0 63962 92 64018
rect 148 63962 216 64018
rect 272 63962 282 64018
rect 0 63894 282 63962
rect 0 63838 92 63894
rect 148 63838 216 63894
rect 272 63838 282 63894
rect 0 63770 282 63838
rect 0 63714 92 63770
rect 148 63714 216 63770
rect 272 63714 282 63770
rect 0 63600 282 63714
rect 81 50600 282 63600
rect 0 50487 282 50600
rect 0 50431 92 50487
rect 148 50431 216 50487
rect 272 50431 282 50487
rect 0 50363 282 50431
rect 0 50307 92 50363
rect 148 50307 216 50363
rect 272 50307 282 50363
rect 0 50239 282 50307
rect 0 50183 92 50239
rect 148 50183 216 50239
rect 272 50183 282 50239
rect 0 50115 282 50183
rect 0 50059 92 50115
rect 148 50059 216 50115
rect 272 50059 282 50115
rect 0 49991 282 50059
rect 0 49935 92 49991
rect 148 49935 216 49991
rect 272 49935 282 49991
rect 0 49867 282 49935
rect 0 49811 92 49867
rect 148 49811 216 49867
rect 272 49811 282 49867
rect 0 49743 282 49811
rect 0 49687 92 49743
rect 148 49687 216 49743
rect 272 49687 282 49743
rect 0 49619 282 49687
rect 0 49563 92 49619
rect 148 49563 216 49619
rect 272 49563 282 49619
rect 0 49495 282 49563
rect 0 49439 92 49495
rect 148 49439 216 49495
rect 272 49439 282 49495
rect 0 49371 282 49439
rect 0 49315 92 49371
rect 148 49315 216 49371
rect 272 49315 282 49371
rect 0 49200 282 49315
rect 81 13611 282 49200
rect 418 68013 604 69054
rect 418 67957 464 68013
rect 520 67957 604 68013
rect 418 67881 604 67957
rect 418 67825 464 67881
rect 520 67825 604 67881
rect 418 67749 604 67825
rect 418 67693 464 67749
rect 520 67693 604 67749
rect 418 67617 604 67693
rect 418 67561 464 67617
rect 520 67561 604 67617
rect 418 67485 604 67561
rect 418 67429 464 67485
rect 520 67429 604 67485
rect 418 67353 604 67429
rect 418 67297 464 67353
rect 520 67297 604 67353
rect 418 67221 604 67297
rect 418 67165 464 67221
rect 520 67165 604 67221
rect 418 67089 604 67165
rect 418 67033 464 67089
rect 520 67033 604 67089
rect 418 66957 604 67033
rect 418 66901 464 66957
rect 520 66901 604 66957
rect 418 60036 604 66901
rect 418 59980 524 60036
rect 580 59980 604 60036
rect 418 59904 604 59980
rect 418 59848 524 59904
rect 580 59848 604 59904
rect 418 59772 604 59848
rect 418 59716 524 59772
rect 580 59716 604 59772
rect 418 59640 604 59716
rect 418 59584 524 59640
rect 580 59584 604 59640
rect 418 59508 604 59584
rect 418 59452 524 59508
rect 580 59452 604 59508
rect 418 59376 604 59452
rect 418 59320 524 59376
rect 580 59320 604 59376
rect 418 59244 604 59320
rect 418 59188 524 59244
rect 580 59188 604 59244
rect 418 59112 604 59188
rect 418 59056 524 59112
rect 580 59056 604 59112
rect 418 58980 604 59056
rect 418 58924 524 58980
rect 580 58924 604 58980
rect 418 56884 604 58924
rect 418 56828 524 56884
rect 580 56828 604 56884
rect 418 56752 604 56828
rect 418 56696 524 56752
rect 580 56696 604 56752
rect 418 56620 604 56696
rect 418 56564 524 56620
rect 580 56564 604 56620
rect 418 56488 604 56564
rect 418 56432 524 56488
rect 580 56432 604 56488
rect 418 56356 604 56432
rect 418 56300 524 56356
rect 580 56300 604 56356
rect 418 56224 604 56300
rect 418 56168 524 56224
rect 580 56168 604 56224
rect 418 56092 604 56168
rect 418 56036 524 56092
rect 580 56036 604 56092
rect 418 55960 604 56036
rect 418 55904 524 55960
rect 580 55904 604 55960
rect 418 55828 604 55904
rect 418 55772 524 55828
rect 580 55772 604 55828
rect 418 55261 604 55772
rect 418 55205 524 55261
rect 580 55205 604 55261
rect 418 55129 604 55205
rect 418 55073 524 55129
rect 580 55073 604 55129
rect 418 54997 604 55073
rect 418 54941 524 54997
rect 580 54941 604 54997
rect 418 54865 604 54941
rect 418 54809 524 54865
rect 580 54809 604 54865
rect 418 54733 604 54809
rect 418 54677 524 54733
rect 580 54677 604 54733
rect 418 54601 604 54677
rect 418 54545 524 54601
rect 580 54545 604 54601
rect 418 54469 604 54545
rect 418 54413 524 54469
rect 580 54413 604 54469
rect 418 54337 604 54413
rect 418 54281 524 54337
rect 580 54281 604 54337
rect 418 54205 604 54281
rect 418 54149 524 54205
rect 580 54149 604 54205
rect 418 53647 604 54149
rect 418 53591 524 53647
rect 580 53591 604 53647
rect 418 53515 604 53591
rect 418 53459 524 53515
rect 580 53459 604 53515
rect 418 53383 604 53459
rect 418 53327 524 53383
rect 580 53327 604 53383
rect 418 53251 604 53327
rect 418 53195 524 53251
rect 580 53195 604 53251
rect 418 53119 604 53195
rect 418 53063 524 53119
rect 580 53063 604 53119
rect 418 52987 604 53063
rect 418 52931 524 52987
rect 580 52931 604 52987
rect 418 52855 604 52931
rect 418 52799 524 52855
rect 580 52799 604 52855
rect 418 52723 604 52799
rect 418 52667 524 52723
rect 580 52667 604 52723
rect 418 52591 604 52667
rect 418 52535 524 52591
rect 580 52535 604 52591
rect 418 45541 604 52535
rect 418 45485 524 45541
rect 580 45485 604 45541
rect 418 45409 604 45485
rect 418 45353 524 45409
rect 580 45353 604 45409
rect 418 45277 604 45353
rect 418 45221 524 45277
rect 580 45221 604 45277
rect 418 45145 604 45221
rect 418 45089 524 45145
rect 580 45089 604 45145
rect 418 45013 604 45089
rect 418 44957 524 45013
rect 580 44957 604 45013
rect 418 44881 604 44957
rect 418 44825 524 44881
rect 580 44825 604 44881
rect 418 44749 604 44825
rect 418 44693 524 44749
rect 580 44693 604 44749
rect 418 44617 604 44693
rect 418 44561 524 44617
rect 580 44561 604 44617
rect 418 44485 604 44561
rect 418 44429 524 44485
rect 580 44429 604 44485
rect 418 44353 604 44429
rect 418 44297 524 44353
rect 580 44297 604 44353
rect 418 44221 604 44297
rect 418 44165 524 44221
rect 580 44165 604 44221
rect 418 44089 604 44165
rect 418 44033 524 44089
rect 580 44033 604 44089
rect 418 43957 604 44033
rect 418 43901 524 43957
rect 580 43901 604 43957
rect 418 43825 604 43901
rect 418 43769 524 43825
rect 580 43769 604 43825
rect 418 43693 604 43769
rect 418 43637 524 43693
rect 580 43637 604 43693
rect 418 43561 604 43637
rect 418 43505 524 43561
rect 580 43505 604 43561
rect 418 43429 604 43505
rect 418 43373 524 43429
rect 580 43373 604 43429
rect 418 43297 604 43373
rect 418 43241 524 43297
rect 580 43241 604 43297
rect 418 43165 604 43241
rect 418 43109 524 43165
rect 580 43109 604 43165
rect 418 43033 604 43109
rect 418 42977 524 43033
rect 580 42977 604 43033
rect 418 42456 604 42977
rect 418 42400 524 42456
rect 580 42400 604 42456
rect 418 42324 604 42400
rect 418 42268 524 42324
rect 580 42268 604 42324
rect 418 42192 604 42268
rect 418 42136 524 42192
rect 580 42136 604 42192
rect 418 42060 604 42136
rect 418 42004 524 42060
rect 580 42004 604 42060
rect 418 41928 604 42004
rect 418 41872 524 41928
rect 580 41872 604 41928
rect 418 41796 604 41872
rect 418 41740 524 41796
rect 580 41740 604 41796
rect 418 41664 604 41740
rect 418 41608 524 41664
rect 580 41608 604 41664
rect 418 41532 604 41608
rect 418 41476 524 41532
rect 580 41476 604 41532
rect 418 41400 604 41476
rect 418 41344 524 41400
rect 580 41344 604 41400
rect 418 39220 604 41344
rect 418 39164 524 39220
rect 580 39164 604 39220
rect 418 39088 604 39164
rect 418 39032 524 39088
rect 580 39032 604 39088
rect 418 38956 604 39032
rect 418 38900 524 38956
rect 580 38900 604 38956
rect 418 38824 604 38900
rect 418 38768 524 38824
rect 580 38768 604 38824
rect 418 38692 604 38768
rect 418 38636 524 38692
rect 580 38636 604 38692
rect 418 38560 604 38636
rect 418 38504 524 38560
rect 580 38504 604 38560
rect 418 38428 604 38504
rect 418 38372 524 38428
rect 580 38372 604 38428
rect 418 38296 604 38372
rect 418 38240 524 38296
rect 580 38240 604 38296
rect 418 38164 604 38240
rect 418 38108 524 38164
rect 580 38108 604 38164
rect 418 38032 604 38108
rect 418 37976 524 38032
rect 580 37976 604 38032
rect 418 37900 604 37976
rect 418 37844 524 37900
rect 580 37844 604 37900
rect 418 37768 604 37844
rect 418 37712 524 37768
rect 580 37712 604 37768
rect 418 37636 604 37712
rect 418 37580 524 37636
rect 580 37580 604 37636
rect 418 37504 604 37580
rect 418 37448 524 37504
rect 580 37448 604 37504
rect 418 37372 604 37448
rect 418 37316 524 37372
rect 580 37316 604 37372
rect 418 37240 604 37316
rect 418 37184 524 37240
rect 580 37184 604 37240
rect 418 37108 604 37184
rect 418 37052 524 37108
rect 580 37052 604 37108
rect 418 36976 604 37052
rect 418 36920 524 36976
rect 580 36920 604 36976
rect 418 36844 604 36920
rect 418 36788 524 36844
rect 580 36788 604 36844
rect 418 36712 604 36788
rect 418 36656 524 36712
rect 580 36656 604 36712
rect 418 35999 604 36656
rect 418 35943 524 35999
rect 580 35943 604 35999
rect 418 35867 604 35943
rect 418 35811 524 35867
rect 580 35811 604 35867
rect 418 35735 604 35811
rect 418 35679 524 35735
rect 580 35679 604 35735
rect 418 35603 604 35679
rect 418 35547 524 35603
rect 580 35547 604 35603
rect 418 35471 604 35547
rect 418 35415 524 35471
rect 580 35415 604 35471
rect 418 35339 604 35415
rect 418 35283 524 35339
rect 580 35283 604 35339
rect 418 35207 604 35283
rect 418 35151 524 35207
rect 580 35151 604 35207
rect 418 35075 604 35151
rect 418 35019 524 35075
rect 580 35019 604 35075
rect 418 34943 604 35019
rect 418 34887 524 34943
rect 580 34887 604 34943
rect 418 34811 604 34887
rect 418 34755 524 34811
rect 580 34755 604 34811
rect 418 34679 604 34755
rect 418 34623 524 34679
rect 580 34623 604 34679
rect 418 34547 604 34623
rect 418 34491 524 34547
rect 580 34491 604 34547
rect 418 34415 604 34491
rect 418 34359 524 34415
rect 580 34359 604 34415
rect 418 34283 604 34359
rect 418 34227 524 34283
rect 580 34227 604 34283
rect 418 34151 604 34227
rect 418 34095 524 34151
rect 580 34095 604 34151
rect 418 34019 604 34095
rect 418 33963 524 34019
rect 580 33963 604 34019
rect 418 33887 604 33963
rect 418 33831 524 33887
rect 580 33831 604 33887
rect 418 33755 604 33831
rect 418 33699 524 33755
rect 580 33699 604 33755
rect 418 33623 604 33699
rect 418 33567 524 33623
rect 580 33567 604 33623
rect 418 33491 604 33567
rect 418 33435 524 33491
rect 580 33435 604 33491
rect 418 32774 604 33435
rect 418 32718 524 32774
rect 580 32718 604 32774
rect 418 32642 604 32718
rect 418 32586 524 32642
rect 580 32586 604 32642
rect 418 32510 604 32586
rect 418 32454 524 32510
rect 580 32454 604 32510
rect 418 32378 604 32454
rect 418 32322 524 32378
rect 580 32322 604 32378
rect 418 32246 604 32322
rect 418 32190 524 32246
rect 580 32190 604 32246
rect 418 32114 604 32190
rect 418 32058 524 32114
rect 580 32058 604 32114
rect 418 31982 604 32058
rect 418 31926 524 31982
rect 580 31926 604 31982
rect 418 31850 604 31926
rect 418 31794 524 31850
rect 580 31794 604 31850
rect 418 31718 604 31794
rect 418 31662 524 31718
rect 580 31662 604 31718
rect 418 31586 604 31662
rect 418 31530 524 31586
rect 580 31530 604 31586
rect 418 31454 604 31530
rect 418 31398 524 31454
rect 580 31398 604 31454
rect 418 31322 604 31398
rect 418 31266 524 31322
rect 580 31266 604 31322
rect 418 31190 604 31266
rect 418 31134 524 31190
rect 580 31134 604 31190
rect 418 31058 604 31134
rect 418 31002 524 31058
rect 580 31002 604 31058
rect 418 30926 604 31002
rect 418 30870 524 30926
rect 580 30870 604 30926
rect 418 30794 604 30870
rect 418 30738 524 30794
rect 580 30738 604 30794
rect 418 30662 604 30738
rect 418 30606 524 30662
rect 580 30606 604 30662
rect 418 30530 604 30606
rect 418 30474 524 30530
rect 580 30474 604 30530
rect 418 30398 604 30474
rect 418 30342 524 30398
rect 580 30342 604 30398
rect 418 30266 604 30342
rect 418 30210 524 30266
rect 580 30210 604 30266
rect 418 29632 604 30210
rect 418 29576 524 29632
rect 580 29576 604 29632
rect 418 29500 604 29576
rect 418 29444 524 29500
rect 580 29444 604 29500
rect 418 29368 604 29444
rect 418 29312 524 29368
rect 580 29312 604 29368
rect 418 29236 604 29312
rect 418 29180 524 29236
rect 580 29180 604 29236
rect 418 29104 604 29180
rect 418 29048 524 29104
rect 580 29048 604 29104
rect 418 28972 604 29048
rect 418 28916 524 28972
rect 580 28916 604 28972
rect 418 28840 604 28916
rect 418 28784 524 28840
rect 580 28784 604 28840
rect 418 28708 604 28784
rect 418 28652 524 28708
rect 580 28652 604 28708
rect 418 28576 604 28652
rect 418 28520 524 28576
rect 580 28520 604 28576
rect 418 28444 604 28520
rect 418 28388 524 28444
rect 580 28388 604 28444
rect 418 28312 604 28388
rect 418 28256 524 28312
rect 580 28256 604 28312
rect 418 28180 604 28256
rect 418 28124 524 28180
rect 580 28124 604 28180
rect 418 28048 604 28124
rect 418 27992 524 28048
rect 580 27992 604 28048
rect 418 27916 604 27992
rect 418 27860 524 27916
rect 580 27860 604 27916
rect 418 27784 604 27860
rect 418 27728 524 27784
rect 580 27728 604 27784
rect 418 27652 604 27728
rect 418 27596 524 27652
rect 580 27596 604 27652
rect 418 27520 604 27596
rect 418 27464 524 27520
rect 580 27464 604 27520
rect 418 27388 604 27464
rect 418 27332 524 27388
rect 580 27332 604 27388
rect 418 27256 604 27332
rect 418 27200 524 27256
rect 580 27200 604 27256
rect 418 27124 604 27200
rect 418 27068 524 27124
rect 580 27068 604 27124
rect 418 24857 604 27068
rect 418 24801 524 24857
rect 580 24801 604 24857
rect 418 24725 604 24801
rect 418 24669 524 24725
rect 580 24669 604 24725
rect 418 24593 604 24669
rect 418 24537 524 24593
rect 580 24537 604 24593
rect 418 24461 604 24537
rect 418 24405 524 24461
rect 580 24405 604 24461
rect 418 24329 604 24405
rect 418 24273 524 24329
rect 580 24273 604 24329
rect 418 24197 604 24273
rect 418 24141 524 24197
rect 580 24141 604 24197
rect 418 24065 604 24141
rect 418 24009 524 24065
rect 580 24009 604 24065
rect 418 23933 604 24009
rect 418 23877 524 23933
rect 580 23877 604 23933
rect 418 23801 604 23877
rect 418 23745 524 23801
rect 580 23745 604 23801
rect 418 23563 604 23745
rect 707 13108 763 69958
rect 922 63321 1130 69075
rect 922 63265 932 63321
rect 988 63265 1064 63321
rect 1120 63265 1130 63321
rect 922 63189 1130 63265
rect 922 63133 932 63189
rect 988 63133 1064 63189
rect 1120 63133 1130 63189
rect 922 63057 1130 63133
rect 922 63001 932 63057
rect 988 63001 1064 63057
rect 1120 63001 1130 63057
rect 922 62925 1130 63001
rect 922 62869 932 62925
rect 988 62869 1064 62925
rect 1120 62869 1130 62925
rect 922 62793 1130 62869
rect 922 62737 932 62793
rect 988 62737 1064 62793
rect 1120 62737 1130 62793
rect 922 62661 1130 62737
rect 922 62605 932 62661
rect 988 62605 1064 62661
rect 1120 62605 1130 62661
rect 922 62529 1130 62605
rect 922 62473 932 62529
rect 988 62473 1064 62529
rect 1120 62473 1130 62529
rect 922 62397 1130 62473
rect 922 62341 932 62397
rect 988 62341 1064 62397
rect 1120 62341 1130 62397
rect 922 62265 1130 62341
rect 922 62209 932 62265
rect 988 62209 1064 62265
rect 1120 62209 1130 62265
rect 922 62133 1130 62209
rect 922 62077 932 62133
rect 988 62077 1064 62133
rect 1120 62077 1130 62133
rect 922 62067 1130 62077
rect 921 52139 1129 52149
rect 921 52083 931 52139
rect 987 52083 1063 52139
rect 1119 52083 1129 52139
rect 921 52007 1129 52083
rect 921 51951 931 52007
rect 987 51951 1063 52007
rect 1119 51951 1129 52007
rect 921 51875 1129 51951
rect 921 51819 931 51875
rect 987 51819 1063 51875
rect 1119 51819 1129 51875
rect 921 51743 1129 51819
rect 921 51687 931 51743
rect 987 51687 1063 51743
rect 1119 51687 1129 51743
rect 921 51611 1129 51687
rect 921 51555 931 51611
rect 987 51555 1063 51611
rect 1119 51555 1129 51611
rect 921 51479 1129 51555
rect 921 51423 931 51479
rect 987 51423 1063 51479
rect 1119 51423 1129 51479
rect 921 51347 1129 51423
rect 921 51291 931 51347
rect 987 51291 1063 51347
rect 1119 51291 1129 51347
rect 921 51215 1129 51291
rect 921 51159 931 51215
rect 987 51159 1063 51215
rect 1119 51159 1129 51215
rect 921 51083 1129 51159
rect 921 51027 931 51083
rect 987 51027 1063 51083
rect 1119 51027 1129 51083
rect 921 50951 1129 51027
rect 921 50895 931 50951
rect 987 50895 1063 50951
rect 1119 50895 1129 50951
rect 921 50885 1129 50895
rect 1290 13108 1346 69958
rect 1426 69610 1591 69629
rect 1426 69554 1507 69610
rect 1563 69554 1591 69610
rect 1426 69478 1591 69554
rect 1426 69422 1507 69478
rect 1563 69422 1591 69478
rect 1426 69346 1591 69422
rect 1426 69290 1507 69346
rect 1563 69290 1591 69346
rect 1426 69214 1591 69290
rect 1426 69158 1507 69214
rect 1563 69158 1591 69214
rect 1426 69082 1591 69158
rect 1426 69026 1507 69082
rect 1563 69026 1591 69082
rect 1426 68950 1591 69026
rect 1426 68894 1507 68950
rect 1563 68894 1591 68950
rect 1426 68818 1591 68894
rect 1426 68762 1507 68818
rect 1563 68762 1591 68818
rect 1426 68686 1591 68762
rect 1426 68630 1507 68686
rect 1563 68630 1591 68686
rect 1426 68554 1591 68630
rect 1426 68498 1507 68554
rect 1563 68498 1591 68554
rect 1426 66473 1591 68498
rect 1426 66417 1447 66473
rect 1503 66417 1591 66473
rect 1426 66341 1591 66417
rect 1426 66285 1447 66341
rect 1503 66285 1591 66341
rect 1426 66209 1591 66285
rect 1426 66153 1447 66209
rect 1503 66153 1591 66209
rect 1426 66077 1591 66153
rect 1426 66021 1447 66077
rect 1503 66021 1591 66077
rect 1426 65945 1591 66021
rect 1426 65889 1447 65945
rect 1503 65889 1591 65945
rect 1426 65813 1591 65889
rect 1426 65757 1447 65813
rect 1503 65757 1591 65813
rect 1426 65681 1591 65757
rect 1426 65625 1447 65681
rect 1503 65625 1591 65681
rect 1426 65549 1591 65625
rect 1426 65493 1447 65549
rect 1503 65493 1591 65549
rect 1426 65417 1591 65493
rect 1426 65361 1447 65417
rect 1503 65361 1591 65417
rect 1426 61677 1591 65361
rect 1426 61621 1447 61677
rect 1503 61621 1591 61677
rect 1426 61545 1591 61621
rect 1426 61489 1447 61545
rect 1503 61489 1591 61545
rect 1426 61413 1591 61489
rect 1426 61357 1447 61413
rect 1503 61357 1591 61413
rect 1426 61281 1591 61357
rect 1426 61225 1447 61281
rect 1503 61225 1591 61281
rect 1426 61149 1591 61225
rect 1426 61093 1447 61149
rect 1503 61093 1591 61149
rect 1426 61017 1591 61093
rect 1426 60961 1447 61017
rect 1503 60961 1591 61017
rect 1426 60885 1591 60961
rect 1426 60829 1447 60885
rect 1503 60829 1591 60885
rect 1426 60753 1591 60829
rect 1426 60697 1447 60753
rect 1503 60697 1591 60753
rect 1426 60621 1591 60697
rect 1426 60565 1447 60621
rect 1503 60565 1591 60621
rect 1426 58439 1591 60565
rect 1426 58383 1447 58439
rect 1503 58383 1591 58439
rect 1426 58307 1591 58383
rect 1426 58251 1447 58307
rect 1503 58251 1591 58307
rect 1426 58175 1591 58251
rect 1426 58119 1447 58175
rect 1503 58119 1591 58175
rect 1426 58043 1591 58119
rect 1426 57987 1447 58043
rect 1503 57987 1591 58043
rect 1426 57911 1591 57987
rect 1426 57855 1447 57911
rect 1503 57855 1591 57911
rect 1426 57779 1591 57855
rect 1426 57723 1447 57779
rect 1503 57723 1591 57779
rect 1426 57647 1591 57723
rect 1426 57591 1447 57647
rect 1503 57591 1591 57647
rect 1426 57515 1591 57591
rect 1426 57459 1447 57515
rect 1503 57459 1591 57515
rect 1426 57383 1591 57459
rect 1426 57327 1447 57383
rect 1503 57327 1591 57383
rect 1426 48765 1591 57327
rect 1426 48709 1447 48765
rect 1503 48709 1591 48765
rect 1426 48633 1591 48709
rect 1426 48577 1447 48633
rect 1503 48577 1591 48633
rect 1426 48501 1591 48577
rect 1426 48445 1447 48501
rect 1503 48445 1591 48501
rect 1426 48369 1591 48445
rect 1426 48313 1447 48369
rect 1503 48313 1591 48369
rect 1426 48237 1591 48313
rect 1426 48181 1447 48237
rect 1503 48181 1591 48237
rect 1426 48105 1591 48181
rect 1426 48049 1447 48105
rect 1503 48049 1591 48105
rect 1426 47973 1591 48049
rect 1426 47917 1447 47973
rect 1503 47917 1591 47973
rect 1426 47841 1591 47917
rect 1426 47785 1447 47841
rect 1503 47785 1591 47841
rect 1426 47709 1591 47785
rect 1426 47653 1447 47709
rect 1503 47653 1591 47709
rect 1426 47577 1591 47653
rect 1426 47521 1447 47577
rect 1503 47521 1591 47577
rect 1426 47445 1591 47521
rect 1426 47389 1447 47445
rect 1503 47389 1591 47445
rect 1426 47313 1591 47389
rect 1426 47257 1447 47313
rect 1503 47257 1591 47313
rect 1426 47181 1591 47257
rect 1426 47125 1447 47181
rect 1503 47125 1591 47181
rect 1426 47049 1591 47125
rect 1426 46993 1447 47049
rect 1503 46993 1591 47049
rect 1426 46917 1591 46993
rect 1426 46861 1447 46917
rect 1503 46861 1591 46917
rect 1426 46785 1591 46861
rect 1426 46729 1447 46785
rect 1503 46729 1591 46785
rect 1426 46653 1591 46729
rect 1426 46597 1447 46653
rect 1503 46597 1591 46653
rect 1426 46521 1591 46597
rect 1426 46465 1447 46521
rect 1503 46465 1591 46521
rect 1426 46389 1591 46465
rect 1426 46333 1447 46389
rect 1503 46333 1591 46389
rect 1426 46257 1591 46333
rect 1426 46201 1447 46257
rect 1503 46201 1591 46257
rect 1426 40884 1591 46201
rect 1426 40828 1447 40884
rect 1503 40828 1591 40884
rect 1426 40752 1591 40828
rect 1426 40696 1447 40752
rect 1503 40696 1591 40752
rect 1426 40620 1591 40696
rect 1426 40564 1447 40620
rect 1503 40564 1591 40620
rect 1426 40488 1591 40564
rect 1426 40432 1447 40488
rect 1503 40432 1591 40488
rect 1426 40356 1591 40432
rect 1426 40300 1447 40356
rect 1503 40300 1591 40356
rect 1426 40224 1591 40300
rect 1426 40168 1447 40224
rect 1503 40168 1591 40224
rect 1426 40092 1591 40168
rect 1426 40036 1447 40092
rect 1503 40036 1591 40092
rect 1426 39960 1591 40036
rect 1426 39904 1447 39960
rect 1503 39904 1591 39960
rect 1426 39828 1591 39904
rect 1426 39772 1447 39828
rect 1503 39772 1591 39828
rect 1426 26490 1591 39772
rect 1426 26434 1447 26490
rect 1503 26434 1591 26490
rect 1426 26358 1591 26434
rect 1426 26302 1447 26358
rect 1503 26302 1591 26358
rect 1426 26226 1591 26302
rect 1426 26170 1447 26226
rect 1503 26170 1591 26226
rect 1426 26094 1591 26170
rect 1426 26038 1447 26094
rect 1503 26038 1591 26094
rect 1426 25962 1591 26038
rect 1426 25906 1447 25962
rect 1503 25906 1591 25962
rect 1426 25830 1591 25906
rect 1426 25774 1447 25830
rect 1503 25774 1591 25830
rect 1426 25698 1591 25774
rect 1426 25642 1447 25698
rect 1503 25642 1591 25698
rect 1426 25566 1591 25642
rect 1426 25510 1447 25566
rect 1503 25510 1591 25566
rect 1426 25434 1591 25510
rect 1426 25378 1447 25434
rect 1503 25378 1591 25434
rect 1426 23151 1591 25378
rect 1426 23095 1447 23151
rect 1503 23095 1591 23151
rect 1426 23019 1591 23095
rect 1426 22963 1447 23019
rect 1503 22963 1591 23019
rect 1426 22887 1591 22963
rect 1426 22831 1447 22887
rect 1503 22831 1591 22887
rect 1426 22755 1591 22831
rect 1426 22699 1447 22755
rect 1503 22699 1591 22755
rect 1426 22623 1591 22699
rect 1426 22567 1447 22623
rect 1503 22567 1591 22623
rect 1426 22491 1591 22567
rect 1426 22435 1447 22491
rect 1503 22435 1591 22491
rect 1426 22359 1591 22435
rect 1426 22303 1447 22359
rect 1503 22303 1591 22359
rect 1426 22227 1591 22303
rect 1426 22171 1447 22227
rect 1503 22171 1591 22227
rect 1426 22095 1591 22171
rect 1426 22039 1447 22095
rect 1503 22039 1591 22095
rect 1426 21963 1591 22039
rect 1426 21907 1447 21963
rect 1503 21907 1591 21963
rect 1426 21831 1591 21907
rect 1426 21775 1447 21831
rect 1503 21775 1591 21831
rect 1426 21699 1591 21775
rect 1426 21643 1447 21699
rect 1503 21643 1591 21699
rect 1426 21567 1591 21643
rect 1426 21511 1447 21567
rect 1503 21511 1591 21567
rect 1426 21435 1591 21511
rect 1426 21379 1447 21435
rect 1503 21379 1591 21435
rect 1426 21303 1591 21379
rect 1426 21247 1447 21303
rect 1503 21247 1591 21303
rect 1426 21171 1591 21247
rect 1426 21115 1447 21171
rect 1503 21115 1591 21171
rect 1426 21039 1591 21115
rect 1426 20983 1447 21039
rect 1503 20983 1591 21039
rect 1426 20907 1591 20983
rect 1426 20851 1447 20907
rect 1503 20851 1591 20907
rect 1426 20775 1591 20851
rect 1426 20719 1447 20775
rect 1503 20719 1591 20775
rect 1426 20643 1591 20719
rect 1426 20587 1447 20643
rect 1503 20587 1591 20643
rect 1426 20004 1591 20587
rect 1426 19948 1447 20004
rect 1503 19948 1591 20004
rect 1426 19872 1591 19948
rect 1426 19816 1447 19872
rect 1503 19816 1591 19872
rect 1426 19740 1591 19816
rect 1426 19684 1447 19740
rect 1503 19684 1591 19740
rect 1426 19608 1591 19684
rect 1426 19552 1447 19608
rect 1503 19552 1591 19608
rect 1426 19476 1591 19552
rect 1426 19420 1447 19476
rect 1503 19420 1591 19476
rect 1426 19344 1591 19420
rect 1426 19288 1447 19344
rect 1503 19288 1591 19344
rect 1426 19212 1591 19288
rect 1426 19156 1447 19212
rect 1503 19156 1591 19212
rect 1426 19080 1591 19156
rect 1426 19024 1447 19080
rect 1503 19024 1591 19080
rect 1426 18948 1591 19024
rect 1426 18892 1447 18948
rect 1503 18892 1591 18948
rect 1426 18816 1591 18892
rect 1426 18760 1447 18816
rect 1503 18760 1591 18816
rect 1426 18684 1591 18760
rect 1426 18628 1447 18684
rect 1503 18628 1591 18684
rect 1426 18552 1591 18628
rect 1426 18496 1447 18552
rect 1503 18496 1591 18552
rect 1426 18420 1591 18496
rect 1426 18364 1447 18420
rect 1503 18364 1591 18420
rect 1426 18288 1591 18364
rect 1426 18232 1447 18288
rect 1503 18232 1591 18288
rect 1426 18156 1591 18232
rect 1426 18100 1447 18156
rect 1503 18100 1591 18156
rect 1426 18024 1591 18100
rect 1426 17968 1447 18024
rect 1503 17968 1591 18024
rect 1426 17892 1591 17968
rect 1426 17836 1447 17892
rect 1503 17836 1591 17892
rect 1426 17760 1591 17836
rect 1426 17704 1447 17760
rect 1503 17704 1591 17760
rect 1426 17628 1591 17704
rect 1426 17572 1447 17628
rect 1503 17572 1591 17628
rect 1426 17496 1591 17572
rect 1426 17440 1447 17496
rect 1503 17440 1591 17496
rect 1426 16814 1591 17440
rect 1426 16758 1447 16814
rect 1503 16758 1591 16814
rect 1426 16682 1591 16758
rect 1426 16626 1447 16682
rect 1503 16626 1591 16682
rect 1426 16550 1591 16626
rect 1426 16494 1447 16550
rect 1503 16494 1591 16550
rect 1426 16418 1591 16494
rect 1426 16362 1447 16418
rect 1503 16362 1591 16418
rect 1426 16286 1591 16362
rect 1426 16230 1447 16286
rect 1503 16230 1591 16286
rect 1426 16154 1591 16230
rect 1426 16098 1447 16154
rect 1503 16098 1591 16154
rect 1426 16022 1591 16098
rect 1426 15966 1447 16022
rect 1503 15966 1591 16022
rect 1426 15890 1591 15966
rect 1426 15834 1447 15890
rect 1503 15834 1591 15890
rect 1426 15758 1591 15834
rect 1426 15702 1447 15758
rect 1503 15702 1591 15758
rect 1426 15626 1591 15702
rect 1426 15570 1447 15626
rect 1503 15570 1591 15626
rect 1426 15494 1591 15570
rect 1426 15438 1447 15494
rect 1503 15438 1591 15494
rect 1426 15362 1591 15438
rect 1426 15306 1447 15362
rect 1503 15306 1591 15362
rect 1426 15230 1591 15306
rect 1426 15174 1447 15230
rect 1503 15174 1591 15230
rect 1426 15098 1591 15174
rect 1426 15042 1447 15098
rect 1503 15042 1591 15098
rect 1426 14966 1591 15042
rect 1426 14910 1447 14966
rect 1503 14910 1591 14966
rect 1426 14834 1591 14910
rect 1426 14778 1447 14834
rect 1503 14778 1591 14834
rect 1426 14702 1591 14778
rect 1426 14646 1447 14702
rect 1503 14646 1591 14702
rect 1426 14570 1591 14646
rect 1426 14514 1447 14570
rect 1503 14514 1591 14570
rect 1426 14438 1591 14514
rect 1426 14382 1447 14438
rect 1503 14382 1591 14438
rect 1426 14306 1591 14382
rect 1426 14250 1447 14306
rect 1503 14250 1591 14306
rect 1426 14031 1591 14250
rect 1717 64886 2000 69054
rect 1717 64830 1728 64886
rect 1784 64830 1852 64886
rect 1908 64830 2000 64886
rect 1717 64762 2000 64830
rect 1717 64706 1728 64762
rect 1784 64706 1852 64762
rect 1908 64706 2000 64762
rect 1717 64638 2000 64706
rect 1717 64582 1728 64638
rect 1784 64582 1852 64638
rect 1908 64582 2000 64638
rect 1717 64514 2000 64582
rect 1717 64458 1728 64514
rect 1784 64458 1852 64514
rect 1908 64458 2000 64514
rect 1717 64390 2000 64458
rect 1717 64334 1728 64390
rect 1784 64334 1852 64390
rect 1908 64334 2000 64390
rect 1717 64266 2000 64334
rect 1717 64210 1728 64266
rect 1784 64210 1852 64266
rect 1908 64210 2000 64266
rect 1717 64142 2000 64210
rect 1717 64086 1728 64142
rect 1784 64086 1852 64142
rect 1908 64086 2000 64142
rect 1717 64018 2000 64086
rect 1717 63962 1728 64018
rect 1784 63962 1852 64018
rect 1908 63962 2000 64018
rect 1717 63894 2000 63962
rect 1717 63838 1728 63894
rect 1784 63838 1852 63894
rect 1908 63838 2000 63894
rect 1717 63770 2000 63838
rect 1717 63714 1728 63770
rect 1784 63714 1852 63770
rect 1908 63714 2000 63770
rect 1717 63600 2000 63714
rect 1717 50600 1918 63600
rect 1717 50487 2000 50600
rect 1717 50431 1728 50487
rect 1784 50431 1852 50487
rect 1908 50431 2000 50487
rect 1717 50363 2000 50431
rect 1717 50307 1728 50363
rect 1784 50307 1852 50363
rect 1908 50307 2000 50363
rect 1717 50239 2000 50307
rect 1717 50183 1728 50239
rect 1784 50183 1852 50239
rect 1908 50183 2000 50239
rect 1717 50115 2000 50183
rect 1717 50059 1728 50115
rect 1784 50059 1852 50115
rect 1908 50059 2000 50115
rect 1717 49991 2000 50059
rect 1717 49935 1728 49991
rect 1784 49935 1852 49991
rect 1908 49935 2000 49991
rect 1717 49867 2000 49935
rect 1717 49811 1728 49867
rect 1784 49811 1852 49867
rect 1908 49811 2000 49867
rect 1717 49743 2000 49811
rect 1717 49687 1728 49743
rect 1784 49687 1852 49743
rect 1908 49687 2000 49743
rect 1717 49619 2000 49687
rect 1717 49563 1728 49619
rect 1784 49563 1852 49619
rect 1908 49563 2000 49619
rect 1717 49495 2000 49563
rect 1717 49439 1728 49495
rect 1784 49439 1852 49495
rect 1908 49439 2000 49495
rect 1717 49371 2000 49439
rect 1717 49315 1728 49371
rect 1784 49315 1852 49371
rect 1908 49315 2000 49371
rect 1717 49200 2000 49315
rect 1717 13611 1918 49200
<< via2 >>
rect 92 64884 148 64886
rect 92 64832 94 64884
rect 94 64832 146 64884
rect 146 64832 148 64884
rect 92 64830 148 64832
rect 216 64884 272 64886
rect 216 64832 218 64884
rect 218 64832 270 64884
rect 270 64832 272 64884
rect 216 64830 272 64832
rect 92 64760 148 64762
rect 92 64708 94 64760
rect 94 64708 146 64760
rect 146 64708 148 64760
rect 92 64706 148 64708
rect 216 64760 272 64762
rect 216 64708 218 64760
rect 218 64708 270 64760
rect 270 64708 272 64760
rect 216 64706 272 64708
rect 92 64636 148 64638
rect 92 64584 94 64636
rect 94 64584 146 64636
rect 146 64584 148 64636
rect 92 64582 148 64584
rect 216 64636 272 64638
rect 216 64584 218 64636
rect 218 64584 270 64636
rect 270 64584 272 64636
rect 216 64582 272 64584
rect 92 64512 148 64514
rect 92 64460 94 64512
rect 94 64460 146 64512
rect 146 64460 148 64512
rect 92 64458 148 64460
rect 216 64512 272 64514
rect 216 64460 218 64512
rect 218 64460 270 64512
rect 270 64460 272 64512
rect 216 64458 272 64460
rect 92 64388 148 64390
rect 92 64336 94 64388
rect 94 64336 146 64388
rect 146 64336 148 64388
rect 92 64334 148 64336
rect 216 64388 272 64390
rect 216 64336 218 64388
rect 218 64336 270 64388
rect 270 64336 272 64388
rect 216 64334 272 64336
rect 92 64264 148 64266
rect 92 64212 94 64264
rect 94 64212 146 64264
rect 146 64212 148 64264
rect 92 64210 148 64212
rect 216 64264 272 64266
rect 216 64212 218 64264
rect 218 64212 270 64264
rect 270 64212 272 64264
rect 216 64210 272 64212
rect 92 64140 148 64142
rect 92 64088 94 64140
rect 94 64088 146 64140
rect 146 64088 148 64140
rect 92 64086 148 64088
rect 216 64140 272 64142
rect 216 64088 218 64140
rect 218 64088 270 64140
rect 270 64088 272 64140
rect 216 64086 272 64088
rect 92 64016 148 64018
rect 92 63964 94 64016
rect 94 63964 146 64016
rect 146 63964 148 64016
rect 92 63962 148 63964
rect 216 64016 272 64018
rect 216 63964 218 64016
rect 218 63964 270 64016
rect 270 63964 272 64016
rect 216 63962 272 63964
rect 92 63892 148 63894
rect 92 63840 94 63892
rect 94 63840 146 63892
rect 146 63840 148 63892
rect 92 63838 148 63840
rect 216 63892 272 63894
rect 216 63840 218 63892
rect 218 63840 270 63892
rect 270 63840 272 63892
rect 216 63838 272 63840
rect 92 63768 148 63770
rect 92 63716 94 63768
rect 94 63716 146 63768
rect 146 63716 148 63768
rect 92 63714 148 63716
rect 216 63768 272 63770
rect 216 63716 218 63768
rect 218 63716 270 63768
rect 270 63716 272 63768
rect 216 63714 272 63716
rect 92 50485 148 50487
rect 92 50433 94 50485
rect 94 50433 146 50485
rect 146 50433 148 50485
rect 92 50431 148 50433
rect 216 50485 272 50487
rect 216 50433 218 50485
rect 218 50433 270 50485
rect 270 50433 272 50485
rect 216 50431 272 50433
rect 92 50361 148 50363
rect 92 50309 94 50361
rect 94 50309 146 50361
rect 146 50309 148 50361
rect 92 50307 148 50309
rect 216 50361 272 50363
rect 216 50309 218 50361
rect 218 50309 270 50361
rect 270 50309 272 50361
rect 216 50307 272 50309
rect 92 50237 148 50239
rect 92 50185 94 50237
rect 94 50185 146 50237
rect 146 50185 148 50237
rect 92 50183 148 50185
rect 216 50237 272 50239
rect 216 50185 218 50237
rect 218 50185 270 50237
rect 270 50185 272 50237
rect 216 50183 272 50185
rect 92 50113 148 50115
rect 92 50061 94 50113
rect 94 50061 146 50113
rect 146 50061 148 50113
rect 92 50059 148 50061
rect 216 50113 272 50115
rect 216 50061 218 50113
rect 218 50061 270 50113
rect 270 50061 272 50113
rect 216 50059 272 50061
rect 92 49989 148 49991
rect 92 49937 94 49989
rect 94 49937 146 49989
rect 146 49937 148 49989
rect 92 49935 148 49937
rect 216 49989 272 49991
rect 216 49937 218 49989
rect 218 49937 270 49989
rect 270 49937 272 49989
rect 216 49935 272 49937
rect 92 49865 148 49867
rect 92 49813 94 49865
rect 94 49813 146 49865
rect 146 49813 148 49865
rect 92 49811 148 49813
rect 216 49865 272 49867
rect 216 49813 218 49865
rect 218 49813 270 49865
rect 270 49813 272 49865
rect 216 49811 272 49813
rect 92 49741 148 49743
rect 92 49689 94 49741
rect 94 49689 146 49741
rect 146 49689 148 49741
rect 92 49687 148 49689
rect 216 49741 272 49743
rect 216 49689 218 49741
rect 218 49689 270 49741
rect 270 49689 272 49741
rect 216 49687 272 49689
rect 92 49617 148 49619
rect 92 49565 94 49617
rect 94 49565 146 49617
rect 146 49565 148 49617
rect 92 49563 148 49565
rect 216 49617 272 49619
rect 216 49565 218 49617
rect 218 49565 270 49617
rect 270 49565 272 49617
rect 216 49563 272 49565
rect 92 49493 148 49495
rect 92 49441 94 49493
rect 94 49441 146 49493
rect 146 49441 148 49493
rect 92 49439 148 49441
rect 216 49493 272 49495
rect 216 49441 218 49493
rect 218 49441 270 49493
rect 270 49441 272 49493
rect 216 49439 272 49441
rect 92 49369 148 49371
rect 92 49317 94 49369
rect 94 49317 146 49369
rect 146 49317 148 49369
rect 92 49315 148 49317
rect 216 49369 272 49371
rect 216 49317 218 49369
rect 218 49317 270 49369
rect 270 49317 272 49369
rect 216 49315 272 49317
rect 464 67957 520 68013
rect 464 67825 520 67881
rect 464 67693 520 67749
rect 464 67561 520 67617
rect 464 67429 520 67485
rect 464 67297 520 67353
rect 464 67165 520 67221
rect 464 67033 520 67089
rect 464 66901 520 66957
rect 524 59980 580 60036
rect 524 59848 580 59904
rect 524 59716 580 59772
rect 524 59584 580 59640
rect 524 59452 580 59508
rect 524 59320 580 59376
rect 524 59188 580 59244
rect 524 59056 580 59112
rect 524 58924 580 58980
rect 524 56828 580 56884
rect 524 56696 580 56752
rect 524 56564 580 56620
rect 524 56432 580 56488
rect 524 56300 580 56356
rect 524 56168 580 56224
rect 524 56036 580 56092
rect 524 55904 580 55960
rect 524 55772 580 55828
rect 524 55205 580 55261
rect 524 55073 580 55129
rect 524 54941 580 54997
rect 524 54809 580 54865
rect 524 54677 580 54733
rect 524 54545 580 54601
rect 524 54413 580 54469
rect 524 54281 580 54337
rect 524 54149 580 54205
rect 524 53591 580 53647
rect 524 53459 580 53515
rect 524 53327 580 53383
rect 524 53195 580 53251
rect 524 53063 580 53119
rect 524 52931 580 52987
rect 524 52799 580 52855
rect 524 52667 580 52723
rect 524 52535 580 52591
rect 524 45485 580 45541
rect 524 45353 580 45409
rect 524 45221 580 45277
rect 524 45089 580 45145
rect 524 44957 580 45013
rect 524 44825 580 44881
rect 524 44693 580 44749
rect 524 44561 580 44617
rect 524 44429 580 44485
rect 524 44297 580 44353
rect 524 44165 580 44221
rect 524 44033 580 44089
rect 524 43901 580 43957
rect 524 43769 580 43825
rect 524 43637 580 43693
rect 524 43505 580 43561
rect 524 43373 580 43429
rect 524 43241 580 43297
rect 524 43109 580 43165
rect 524 42977 580 43033
rect 524 42400 580 42456
rect 524 42268 580 42324
rect 524 42136 580 42192
rect 524 42004 580 42060
rect 524 41872 580 41928
rect 524 41740 580 41796
rect 524 41608 580 41664
rect 524 41476 580 41532
rect 524 41344 580 41400
rect 524 39164 580 39220
rect 524 39032 580 39088
rect 524 38900 580 38956
rect 524 38768 580 38824
rect 524 38636 580 38692
rect 524 38504 580 38560
rect 524 38372 580 38428
rect 524 38240 580 38296
rect 524 38108 580 38164
rect 524 37976 580 38032
rect 524 37844 580 37900
rect 524 37712 580 37768
rect 524 37580 580 37636
rect 524 37448 580 37504
rect 524 37316 580 37372
rect 524 37184 580 37240
rect 524 37052 580 37108
rect 524 36920 580 36976
rect 524 36788 580 36844
rect 524 36656 580 36712
rect 524 35943 580 35999
rect 524 35811 580 35867
rect 524 35679 580 35735
rect 524 35547 580 35603
rect 524 35415 580 35471
rect 524 35283 580 35339
rect 524 35151 580 35207
rect 524 35019 580 35075
rect 524 34887 580 34943
rect 524 34755 580 34811
rect 524 34623 580 34679
rect 524 34491 580 34547
rect 524 34359 580 34415
rect 524 34227 580 34283
rect 524 34095 580 34151
rect 524 33963 580 34019
rect 524 33831 580 33887
rect 524 33699 580 33755
rect 524 33567 580 33623
rect 524 33435 580 33491
rect 524 32718 580 32774
rect 524 32586 580 32642
rect 524 32454 580 32510
rect 524 32322 580 32378
rect 524 32190 580 32246
rect 524 32058 580 32114
rect 524 31926 580 31982
rect 524 31794 580 31850
rect 524 31662 580 31718
rect 524 31530 580 31586
rect 524 31398 580 31454
rect 524 31266 580 31322
rect 524 31134 580 31190
rect 524 31002 580 31058
rect 524 30870 580 30926
rect 524 30738 580 30794
rect 524 30606 580 30662
rect 524 30474 580 30530
rect 524 30342 580 30398
rect 524 30210 580 30266
rect 524 29576 580 29632
rect 524 29444 580 29500
rect 524 29312 580 29368
rect 524 29180 580 29236
rect 524 29048 580 29104
rect 524 28916 580 28972
rect 524 28784 580 28840
rect 524 28652 580 28708
rect 524 28520 580 28576
rect 524 28388 580 28444
rect 524 28256 580 28312
rect 524 28124 580 28180
rect 524 27992 580 28048
rect 524 27860 580 27916
rect 524 27728 580 27784
rect 524 27596 580 27652
rect 524 27464 580 27520
rect 524 27332 580 27388
rect 524 27200 580 27256
rect 524 27068 580 27124
rect 524 24801 580 24857
rect 524 24669 580 24725
rect 524 24537 580 24593
rect 524 24405 580 24461
rect 524 24273 580 24329
rect 524 24141 580 24197
rect 524 24009 580 24065
rect 524 23877 580 23933
rect 524 23745 580 23801
rect 932 63265 988 63321
rect 1064 63265 1120 63321
rect 932 63133 988 63189
rect 1064 63133 1120 63189
rect 932 63001 988 63057
rect 1064 63001 1120 63057
rect 932 62869 988 62925
rect 1064 62869 1120 62925
rect 932 62737 988 62793
rect 1064 62737 1120 62793
rect 932 62605 988 62661
rect 1064 62605 1120 62661
rect 932 62473 988 62529
rect 1064 62473 1120 62529
rect 932 62341 988 62397
rect 1064 62341 1120 62397
rect 932 62209 988 62265
rect 1064 62209 1120 62265
rect 932 62077 988 62133
rect 1064 62077 1120 62133
rect 931 52083 987 52139
rect 1063 52083 1119 52139
rect 931 51951 987 52007
rect 1063 51951 1119 52007
rect 931 51819 987 51875
rect 1063 51819 1119 51875
rect 931 51687 987 51743
rect 1063 51687 1119 51743
rect 931 51555 987 51611
rect 1063 51555 1119 51611
rect 931 51423 987 51479
rect 1063 51423 1119 51479
rect 931 51291 987 51347
rect 1063 51291 1119 51347
rect 931 51159 987 51215
rect 1063 51159 1119 51215
rect 931 51027 987 51083
rect 1063 51027 1119 51083
rect 931 50895 987 50951
rect 1063 50895 1119 50951
rect 1507 69554 1563 69610
rect 1507 69422 1563 69478
rect 1507 69290 1563 69346
rect 1507 69158 1563 69214
rect 1507 69026 1563 69082
rect 1507 68894 1563 68950
rect 1507 68762 1563 68818
rect 1507 68630 1563 68686
rect 1507 68498 1563 68554
rect 1447 66417 1503 66473
rect 1447 66285 1503 66341
rect 1447 66153 1503 66209
rect 1447 66021 1503 66077
rect 1447 65889 1503 65945
rect 1447 65757 1503 65813
rect 1447 65625 1503 65681
rect 1447 65493 1503 65549
rect 1447 65361 1503 65417
rect 1447 61621 1503 61677
rect 1447 61489 1503 61545
rect 1447 61357 1503 61413
rect 1447 61225 1503 61281
rect 1447 61093 1503 61149
rect 1447 60961 1503 61017
rect 1447 60829 1503 60885
rect 1447 60697 1503 60753
rect 1447 60565 1503 60621
rect 1447 58383 1503 58439
rect 1447 58251 1503 58307
rect 1447 58119 1503 58175
rect 1447 57987 1503 58043
rect 1447 57855 1503 57911
rect 1447 57723 1503 57779
rect 1447 57591 1503 57647
rect 1447 57459 1503 57515
rect 1447 57327 1503 57383
rect 1447 48709 1503 48765
rect 1447 48577 1503 48633
rect 1447 48445 1503 48501
rect 1447 48313 1503 48369
rect 1447 48181 1503 48237
rect 1447 48049 1503 48105
rect 1447 47917 1503 47973
rect 1447 47785 1503 47841
rect 1447 47653 1503 47709
rect 1447 47521 1503 47577
rect 1447 47389 1503 47445
rect 1447 47257 1503 47313
rect 1447 47125 1503 47181
rect 1447 46993 1503 47049
rect 1447 46861 1503 46917
rect 1447 46729 1503 46785
rect 1447 46597 1503 46653
rect 1447 46465 1503 46521
rect 1447 46333 1503 46389
rect 1447 46201 1503 46257
rect 1447 40828 1503 40884
rect 1447 40696 1503 40752
rect 1447 40564 1503 40620
rect 1447 40432 1503 40488
rect 1447 40300 1503 40356
rect 1447 40168 1503 40224
rect 1447 40036 1503 40092
rect 1447 39904 1503 39960
rect 1447 39772 1503 39828
rect 1447 26434 1503 26490
rect 1447 26302 1503 26358
rect 1447 26170 1503 26226
rect 1447 26038 1503 26094
rect 1447 25906 1503 25962
rect 1447 25774 1503 25830
rect 1447 25642 1503 25698
rect 1447 25510 1503 25566
rect 1447 25378 1503 25434
rect 1447 23095 1503 23151
rect 1447 22963 1503 23019
rect 1447 22831 1503 22887
rect 1447 22699 1503 22755
rect 1447 22567 1503 22623
rect 1447 22435 1503 22491
rect 1447 22303 1503 22359
rect 1447 22171 1503 22227
rect 1447 22039 1503 22095
rect 1447 21907 1503 21963
rect 1447 21775 1503 21831
rect 1447 21643 1503 21699
rect 1447 21511 1503 21567
rect 1447 21379 1503 21435
rect 1447 21247 1503 21303
rect 1447 21115 1503 21171
rect 1447 20983 1503 21039
rect 1447 20851 1503 20907
rect 1447 20719 1503 20775
rect 1447 20587 1503 20643
rect 1447 19948 1503 20004
rect 1447 19816 1503 19872
rect 1447 19684 1503 19740
rect 1447 19552 1503 19608
rect 1447 19420 1503 19476
rect 1447 19288 1503 19344
rect 1447 19156 1503 19212
rect 1447 19024 1503 19080
rect 1447 18892 1503 18948
rect 1447 18760 1503 18816
rect 1447 18628 1503 18684
rect 1447 18496 1503 18552
rect 1447 18364 1503 18420
rect 1447 18232 1503 18288
rect 1447 18100 1503 18156
rect 1447 17968 1503 18024
rect 1447 17836 1503 17892
rect 1447 17704 1503 17760
rect 1447 17572 1503 17628
rect 1447 17440 1503 17496
rect 1447 16758 1503 16814
rect 1447 16626 1503 16682
rect 1447 16494 1503 16550
rect 1447 16362 1503 16418
rect 1447 16230 1503 16286
rect 1447 16098 1503 16154
rect 1447 15966 1503 16022
rect 1447 15834 1503 15890
rect 1447 15702 1503 15758
rect 1447 15570 1503 15626
rect 1447 15438 1503 15494
rect 1447 15306 1503 15362
rect 1447 15174 1503 15230
rect 1447 15042 1503 15098
rect 1447 14910 1503 14966
rect 1447 14778 1503 14834
rect 1447 14646 1503 14702
rect 1447 14514 1503 14570
rect 1447 14382 1503 14438
rect 1447 14250 1503 14306
rect 1728 64884 1784 64886
rect 1728 64832 1730 64884
rect 1730 64832 1782 64884
rect 1782 64832 1784 64884
rect 1728 64830 1784 64832
rect 1852 64884 1908 64886
rect 1852 64832 1854 64884
rect 1854 64832 1906 64884
rect 1906 64832 1908 64884
rect 1852 64830 1908 64832
rect 1728 64760 1784 64762
rect 1728 64708 1730 64760
rect 1730 64708 1782 64760
rect 1782 64708 1784 64760
rect 1728 64706 1784 64708
rect 1852 64760 1908 64762
rect 1852 64708 1854 64760
rect 1854 64708 1906 64760
rect 1906 64708 1908 64760
rect 1852 64706 1908 64708
rect 1728 64636 1784 64638
rect 1728 64584 1730 64636
rect 1730 64584 1782 64636
rect 1782 64584 1784 64636
rect 1728 64582 1784 64584
rect 1852 64636 1908 64638
rect 1852 64584 1854 64636
rect 1854 64584 1906 64636
rect 1906 64584 1908 64636
rect 1852 64582 1908 64584
rect 1728 64512 1784 64514
rect 1728 64460 1730 64512
rect 1730 64460 1782 64512
rect 1782 64460 1784 64512
rect 1728 64458 1784 64460
rect 1852 64512 1908 64514
rect 1852 64460 1854 64512
rect 1854 64460 1906 64512
rect 1906 64460 1908 64512
rect 1852 64458 1908 64460
rect 1728 64388 1784 64390
rect 1728 64336 1730 64388
rect 1730 64336 1782 64388
rect 1782 64336 1784 64388
rect 1728 64334 1784 64336
rect 1852 64388 1908 64390
rect 1852 64336 1854 64388
rect 1854 64336 1906 64388
rect 1906 64336 1908 64388
rect 1852 64334 1908 64336
rect 1728 64264 1784 64266
rect 1728 64212 1730 64264
rect 1730 64212 1782 64264
rect 1782 64212 1784 64264
rect 1728 64210 1784 64212
rect 1852 64264 1908 64266
rect 1852 64212 1854 64264
rect 1854 64212 1906 64264
rect 1906 64212 1908 64264
rect 1852 64210 1908 64212
rect 1728 64140 1784 64142
rect 1728 64088 1730 64140
rect 1730 64088 1782 64140
rect 1782 64088 1784 64140
rect 1728 64086 1784 64088
rect 1852 64140 1908 64142
rect 1852 64088 1854 64140
rect 1854 64088 1906 64140
rect 1906 64088 1908 64140
rect 1852 64086 1908 64088
rect 1728 64016 1784 64018
rect 1728 63964 1730 64016
rect 1730 63964 1782 64016
rect 1782 63964 1784 64016
rect 1728 63962 1784 63964
rect 1852 64016 1908 64018
rect 1852 63964 1854 64016
rect 1854 63964 1906 64016
rect 1906 63964 1908 64016
rect 1852 63962 1908 63964
rect 1728 63892 1784 63894
rect 1728 63840 1730 63892
rect 1730 63840 1782 63892
rect 1782 63840 1784 63892
rect 1728 63838 1784 63840
rect 1852 63892 1908 63894
rect 1852 63840 1854 63892
rect 1854 63840 1906 63892
rect 1906 63840 1908 63892
rect 1852 63838 1908 63840
rect 1728 63768 1784 63770
rect 1728 63716 1730 63768
rect 1730 63716 1782 63768
rect 1782 63716 1784 63768
rect 1728 63714 1784 63716
rect 1852 63768 1908 63770
rect 1852 63716 1854 63768
rect 1854 63716 1906 63768
rect 1906 63716 1908 63768
rect 1852 63714 1908 63716
rect 1728 50485 1784 50487
rect 1728 50433 1730 50485
rect 1730 50433 1782 50485
rect 1782 50433 1784 50485
rect 1728 50431 1784 50433
rect 1852 50485 1908 50487
rect 1852 50433 1854 50485
rect 1854 50433 1906 50485
rect 1906 50433 1908 50485
rect 1852 50431 1908 50433
rect 1728 50361 1784 50363
rect 1728 50309 1730 50361
rect 1730 50309 1782 50361
rect 1782 50309 1784 50361
rect 1728 50307 1784 50309
rect 1852 50361 1908 50363
rect 1852 50309 1854 50361
rect 1854 50309 1906 50361
rect 1906 50309 1908 50361
rect 1852 50307 1908 50309
rect 1728 50237 1784 50239
rect 1728 50185 1730 50237
rect 1730 50185 1782 50237
rect 1782 50185 1784 50237
rect 1728 50183 1784 50185
rect 1852 50237 1908 50239
rect 1852 50185 1854 50237
rect 1854 50185 1906 50237
rect 1906 50185 1908 50237
rect 1852 50183 1908 50185
rect 1728 50113 1784 50115
rect 1728 50061 1730 50113
rect 1730 50061 1782 50113
rect 1782 50061 1784 50113
rect 1728 50059 1784 50061
rect 1852 50113 1908 50115
rect 1852 50061 1854 50113
rect 1854 50061 1906 50113
rect 1906 50061 1908 50113
rect 1852 50059 1908 50061
rect 1728 49989 1784 49991
rect 1728 49937 1730 49989
rect 1730 49937 1782 49989
rect 1782 49937 1784 49989
rect 1728 49935 1784 49937
rect 1852 49989 1908 49991
rect 1852 49937 1854 49989
rect 1854 49937 1906 49989
rect 1906 49937 1908 49989
rect 1852 49935 1908 49937
rect 1728 49865 1784 49867
rect 1728 49813 1730 49865
rect 1730 49813 1782 49865
rect 1782 49813 1784 49865
rect 1728 49811 1784 49813
rect 1852 49865 1908 49867
rect 1852 49813 1854 49865
rect 1854 49813 1906 49865
rect 1906 49813 1908 49865
rect 1852 49811 1908 49813
rect 1728 49741 1784 49743
rect 1728 49689 1730 49741
rect 1730 49689 1782 49741
rect 1782 49689 1784 49741
rect 1728 49687 1784 49689
rect 1852 49741 1908 49743
rect 1852 49689 1854 49741
rect 1854 49689 1906 49741
rect 1906 49689 1908 49741
rect 1852 49687 1908 49689
rect 1728 49617 1784 49619
rect 1728 49565 1730 49617
rect 1730 49565 1782 49617
rect 1782 49565 1784 49617
rect 1728 49563 1784 49565
rect 1852 49617 1908 49619
rect 1852 49565 1854 49617
rect 1854 49565 1906 49617
rect 1906 49565 1908 49617
rect 1852 49563 1908 49565
rect 1728 49493 1784 49495
rect 1728 49441 1730 49493
rect 1730 49441 1782 49493
rect 1782 49441 1784 49493
rect 1728 49439 1784 49441
rect 1852 49493 1908 49495
rect 1852 49441 1854 49493
rect 1854 49441 1906 49493
rect 1906 49441 1908 49493
rect 1852 49439 1908 49441
rect 1728 49369 1784 49371
rect 1728 49317 1730 49369
rect 1730 49317 1782 49369
rect 1782 49317 1784 49369
rect 1728 49315 1784 49317
rect 1852 49369 1908 49371
rect 1852 49317 1854 49369
rect 1854 49317 1906 49369
rect 1906 49317 1908 49369
rect 1852 49315 1908 49317
<< metal3 >>
rect 0 69610 2000 69678
rect 0 69554 1507 69610
rect 1563 69554 2000 69610
rect 0 69478 2000 69554
rect 0 69422 1507 69478
rect 1563 69422 2000 69478
rect 0 69346 2000 69422
rect 0 69290 1507 69346
rect 1563 69290 2000 69346
rect 0 69214 2000 69290
rect 0 69158 1507 69214
rect 1563 69158 2000 69214
rect 0 69082 2000 69158
rect 0 69026 1507 69082
rect 1563 69026 2000 69082
rect 0 68950 2000 69026
rect 0 68894 1507 68950
rect 1563 68894 2000 68950
rect 0 68818 2000 68894
rect 0 68762 1507 68818
rect 1563 68762 2000 68818
rect 0 68686 2000 68762
rect 0 68630 1507 68686
rect 1563 68630 2000 68686
rect 0 68554 2000 68630
rect 0 68498 1507 68554
rect 1563 68498 2000 68554
rect 0 68400 2000 68498
rect 0 68013 2000 68200
rect 0 67957 464 68013
rect 520 67957 2000 68013
rect 0 67881 2000 67957
rect 0 67825 464 67881
rect 520 67825 2000 67881
rect 0 67749 2000 67825
rect 0 67693 464 67749
rect 520 67693 2000 67749
rect 0 67617 2000 67693
rect 0 67561 464 67617
rect 520 67561 2000 67617
rect 0 67485 2000 67561
rect 0 67429 464 67485
rect 520 67429 2000 67485
rect 0 67353 2000 67429
rect 0 67297 464 67353
rect 520 67297 2000 67353
rect 0 67221 2000 67297
rect 0 67165 464 67221
rect 520 67165 2000 67221
rect 0 67089 2000 67165
rect 0 67033 464 67089
rect 520 67033 2000 67089
rect 0 66957 2000 67033
rect 0 66901 464 66957
rect 520 66901 2000 66957
rect 0 66800 2000 66901
rect 0 66473 2000 66600
rect 0 66417 1447 66473
rect 1503 66417 2000 66473
rect 0 66341 2000 66417
rect 0 66285 1447 66341
rect 1503 66285 2000 66341
rect 0 66209 2000 66285
rect 0 66153 1447 66209
rect 1503 66153 2000 66209
rect 0 66077 2000 66153
rect 0 66021 1447 66077
rect 1503 66021 2000 66077
rect 0 65945 2000 66021
rect 0 65889 1447 65945
rect 1503 65889 2000 65945
rect 0 65813 2000 65889
rect 0 65757 1447 65813
rect 1503 65757 2000 65813
rect 0 65681 2000 65757
rect 0 65625 1447 65681
rect 1503 65625 2000 65681
rect 0 65549 2000 65625
rect 0 65493 1447 65549
rect 1503 65493 2000 65549
rect 0 65417 2000 65493
rect 0 65361 1447 65417
rect 1503 65361 2000 65417
rect 0 65200 2000 65361
rect 0 64886 2000 65000
rect 0 64830 92 64886
rect 148 64830 216 64886
rect 272 64830 1728 64886
rect 1784 64830 1852 64886
rect 1908 64830 2000 64886
rect 0 64762 2000 64830
rect 0 64706 92 64762
rect 148 64706 216 64762
rect 272 64706 1728 64762
rect 1784 64706 1852 64762
rect 1908 64706 2000 64762
rect 0 64638 2000 64706
rect 0 64582 92 64638
rect 148 64582 216 64638
rect 272 64582 1728 64638
rect 1784 64582 1852 64638
rect 1908 64582 2000 64638
rect 0 64514 2000 64582
rect 0 64458 92 64514
rect 148 64458 216 64514
rect 272 64458 1728 64514
rect 1784 64458 1852 64514
rect 1908 64458 2000 64514
rect 0 64390 2000 64458
rect 0 64334 92 64390
rect 148 64334 216 64390
rect 272 64334 1728 64390
rect 1784 64334 1852 64390
rect 1908 64334 2000 64390
rect 0 64266 2000 64334
rect 0 64210 92 64266
rect 148 64210 216 64266
rect 272 64210 1728 64266
rect 1784 64210 1852 64266
rect 1908 64210 2000 64266
rect 0 64142 2000 64210
rect 0 64086 92 64142
rect 148 64086 216 64142
rect 272 64086 1728 64142
rect 1784 64086 1852 64142
rect 1908 64086 2000 64142
rect 0 64018 2000 64086
rect 0 63962 92 64018
rect 148 63962 216 64018
rect 272 63962 1728 64018
rect 1784 63962 1852 64018
rect 1908 63962 2000 64018
rect 0 63894 2000 63962
rect 0 63838 92 63894
rect 148 63838 216 63894
rect 272 63838 1728 63894
rect 1784 63838 1852 63894
rect 1908 63838 2000 63894
rect 0 63770 2000 63838
rect 0 63714 92 63770
rect 148 63714 216 63770
rect 272 63714 1728 63770
rect 1784 63714 1852 63770
rect 1908 63714 2000 63770
rect 0 63600 2000 63714
rect 0 63321 2000 63400
rect 0 63265 932 63321
rect 988 63265 1064 63321
rect 1120 63265 2000 63321
rect 0 63189 2000 63265
rect 0 63133 932 63189
rect 988 63133 1064 63189
rect 1120 63133 2000 63189
rect 0 63057 2000 63133
rect 0 63001 932 63057
rect 988 63001 1064 63057
rect 1120 63001 2000 63057
rect 0 62925 2000 63001
rect 0 62869 932 62925
rect 988 62869 1064 62925
rect 1120 62869 2000 62925
rect 0 62793 2000 62869
rect 0 62737 932 62793
rect 988 62737 1064 62793
rect 1120 62737 2000 62793
rect 0 62661 2000 62737
rect 0 62605 932 62661
rect 988 62605 1064 62661
rect 1120 62605 2000 62661
rect 0 62529 2000 62605
rect 0 62473 932 62529
rect 988 62473 1064 62529
rect 1120 62473 2000 62529
rect 0 62397 2000 62473
rect 0 62341 932 62397
rect 988 62341 1064 62397
rect 1120 62341 2000 62397
rect 0 62265 2000 62341
rect 0 62209 932 62265
rect 988 62209 1064 62265
rect 1120 62209 2000 62265
rect 0 62133 2000 62209
rect 0 62077 932 62133
rect 988 62077 1064 62133
rect 1120 62077 2000 62133
rect 0 62000 2000 62077
rect 0 61677 2000 61800
rect 0 61621 1447 61677
rect 1503 61621 2000 61677
rect 0 61545 2000 61621
rect 0 61489 1447 61545
rect 1503 61489 2000 61545
rect 0 61413 2000 61489
rect 0 61357 1447 61413
rect 1503 61357 2000 61413
rect 0 61281 2000 61357
rect 0 61225 1447 61281
rect 1503 61225 2000 61281
rect 0 61149 2000 61225
rect 0 61093 1447 61149
rect 1503 61093 2000 61149
rect 0 61017 2000 61093
rect 0 60961 1447 61017
rect 1503 60961 2000 61017
rect 0 60885 2000 60961
rect 0 60829 1447 60885
rect 1503 60829 2000 60885
rect 0 60753 2000 60829
rect 0 60697 1447 60753
rect 1503 60697 2000 60753
rect 0 60621 2000 60697
rect 0 60565 1447 60621
rect 1503 60565 2000 60621
rect 0 60400 2000 60565
rect 0 60036 2000 60200
rect 0 59980 524 60036
rect 580 59980 2000 60036
rect 0 59904 2000 59980
rect 0 59848 524 59904
rect 580 59848 2000 59904
rect 0 59772 2000 59848
rect 0 59716 524 59772
rect 580 59716 2000 59772
rect 0 59640 2000 59716
rect 0 59584 524 59640
rect 580 59584 2000 59640
rect 0 59508 2000 59584
rect 0 59452 524 59508
rect 580 59452 2000 59508
rect 0 59376 2000 59452
rect 0 59320 524 59376
rect 580 59320 2000 59376
rect 0 59244 2000 59320
rect 0 59188 524 59244
rect 580 59188 2000 59244
rect 0 59112 2000 59188
rect 0 59056 524 59112
rect 580 59056 2000 59112
rect 0 58980 2000 59056
rect 0 58924 524 58980
rect 580 58924 2000 58980
rect 0 58800 2000 58924
rect 0 58439 2000 58600
rect 0 58383 1447 58439
rect 1503 58383 2000 58439
rect 0 58307 2000 58383
rect 0 58251 1447 58307
rect 1503 58251 2000 58307
rect 0 58175 2000 58251
rect 0 58119 1447 58175
rect 1503 58119 2000 58175
rect 0 58043 2000 58119
rect 0 57987 1447 58043
rect 1503 57987 2000 58043
rect 0 57911 2000 57987
rect 0 57855 1447 57911
rect 1503 57855 2000 57911
rect 0 57779 2000 57855
rect 0 57723 1447 57779
rect 1503 57723 2000 57779
rect 0 57647 2000 57723
rect 0 57591 1447 57647
rect 1503 57591 2000 57647
rect 0 57515 2000 57591
rect 0 57459 1447 57515
rect 1503 57459 2000 57515
rect 0 57383 2000 57459
rect 0 57327 1447 57383
rect 1503 57327 2000 57383
rect 0 57200 2000 57327
rect 0 56884 2000 57000
rect 0 56828 524 56884
rect 580 56828 2000 56884
rect 0 56752 2000 56828
rect 0 56696 524 56752
rect 580 56696 2000 56752
rect 0 56620 2000 56696
rect 0 56564 524 56620
rect 580 56564 2000 56620
rect 0 56488 2000 56564
rect 0 56432 524 56488
rect 580 56432 2000 56488
rect 0 56356 2000 56432
rect 0 56300 524 56356
rect 580 56300 2000 56356
rect 0 56224 2000 56300
rect 0 56168 524 56224
rect 580 56168 2000 56224
rect 0 56092 2000 56168
rect 0 56036 524 56092
rect 580 56036 2000 56092
rect 0 55960 2000 56036
rect 0 55904 524 55960
rect 580 55904 2000 55960
rect 0 55828 2000 55904
rect 0 55772 524 55828
rect 580 55772 2000 55828
rect 0 55600 2000 55772
rect 0 55261 2000 55400
rect 0 55205 524 55261
rect 580 55205 2000 55261
rect 0 55129 2000 55205
rect 0 55073 524 55129
rect 580 55073 2000 55129
rect 0 54997 2000 55073
rect 0 54941 524 54997
rect 580 54941 2000 54997
rect 0 54865 2000 54941
rect 0 54809 524 54865
rect 580 54809 2000 54865
rect 0 54733 2000 54809
rect 0 54677 524 54733
rect 580 54677 2000 54733
rect 0 54601 2000 54677
rect 0 54545 524 54601
rect 580 54545 2000 54601
rect 0 54469 2000 54545
rect 0 54413 524 54469
rect 580 54413 2000 54469
rect 0 54337 2000 54413
rect 0 54281 524 54337
rect 580 54281 2000 54337
rect 0 54205 2000 54281
rect 0 54149 524 54205
rect 580 54149 2000 54205
rect 0 54000 2000 54149
rect 0 53647 2000 53800
rect 0 53591 524 53647
rect 580 53591 2000 53647
rect 0 53515 2000 53591
rect 0 53459 524 53515
rect 580 53459 2000 53515
rect 0 53383 2000 53459
rect 0 53327 524 53383
rect 580 53327 2000 53383
rect 0 53251 2000 53327
rect 0 53195 524 53251
rect 580 53195 2000 53251
rect 0 53119 2000 53195
rect 0 53063 524 53119
rect 580 53063 2000 53119
rect 0 52987 2000 53063
rect 0 52931 524 52987
rect 580 52931 2000 52987
rect 0 52855 2000 52931
rect 0 52799 524 52855
rect 580 52799 2000 52855
rect 0 52723 2000 52799
rect 0 52667 524 52723
rect 580 52667 2000 52723
rect 0 52591 2000 52667
rect 0 52535 524 52591
rect 580 52535 2000 52591
rect 0 52400 2000 52535
rect 0 52139 2000 52200
rect 0 52083 931 52139
rect 987 52083 1063 52139
rect 1119 52083 2000 52139
rect 0 52007 2000 52083
rect 0 51951 931 52007
rect 987 51951 1063 52007
rect 1119 51951 2000 52007
rect 0 51875 2000 51951
rect 0 51819 931 51875
rect 987 51819 1063 51875
rect 1119 51819 2000 51875
rect 0 51743 2000 51819
rect 0 51687 931 51743
rect 987 51687 1063 51743
rect 1119 51687 2000 51743
rect 0 51611 2000 51687
rect 0 51555 931 51611
rect 987 51555 1063 51611
rect 1119 51555 2000 51611
rect 0 51479 2000 51555
rect 0 51423 931 51479
rect 987 51423 1063 51479
rect 1119 51423 2000 51479
rect 0 51347 2000 51423
rect 0 51291 931 51347
rect 987 51291 1063 51347
rect 1119 51291 2000 51347
rect 0 51215 2000 51291
rect 0 51159 931 51215
rect 987 51159 1063 51215
rect 1119 51159 2000 51215
rect 0 51083 2000 51159
rect 0 51027 931 51083
rect 987 51027 1063 51083
rect 1119 51027 2000 51083
rect 0 50951 2000 51027
rect 0 50895 931 50951
rect 987 50895 1063 50951
rect 1119 50895 2000 50951
rect 0 50800 2000 50895
rect 0 50487 2000 50600
rect 0 50431 92 50487
rect 148 50431 216 50487
rect 272 50431 1728 50487
rect 1784 50431 1852 50487
rect 1908 50431 2000 50487
rect 0 50363 2000 50431
rect 0 50307 92 50363
rect 148 50307 216 50363
rect 272 50307 1728 50363
rect 1784 50307 1852 50363
rect 1908 50307 2000 50363
rect 0 50239 2000 50307
rect 0 50183 92 50239
rect 148 50183 216 50239
rect 272 50183 1728 50239
rect 1784 50183 1852 50239
rect 1908 50183 2000 50239
rect 0 50115 2000 50183
rect 0 50059 92 50115
rect 148 50059 216 50115
rect 272 50059 1728 50115
rect 1784 50059 1852 50115
rect 1908 50059 2000 50115
rect 0 49991 2000 50059
rect 0 49935 92 49991
rect 148 49935 216 49991
rect 272 49935 1728 49991
rect 1784 49935 1852 49991
rect 1908 49935 2000 49991
rect 0 49867 2000 49935
rect 0 49811 92 49867
rect 148 49811 216 49867
rect 272 49811 1728 49867
rect 1784 49811 1852 49867
rect 1908 49811 2000 49867
rect 0 49743 2000 49811
rect 0 49687 92 49743
rect 148 49687 216 49743
rect 272 49687 1728 49743
rect 1784 49687 1852 49743
rect 1908 49687 2000 49743
rect 0 49619 2000 49687
rect 0 49563 92 49619
rect 148 49563 216 49619
rect 272 49563 1728 49619
rect 1784 49563 1852 49619
rect 1908 49563 2000 49619
rect 0 49495 2000 49563
rect 0 49439 92 49495
rect 148 49439 216 49495
rect 272 49439 1728 49495
rect 1784 49439 1852 49495
rect 1908 49439 2000 49495
rect 0 49371 2000 49439
rect 0 49315 92 49371
rect 148 49315 216 49371
rect 272 49315 1728 49371
rect 1784 49315 1852 49371
rect 1908 49315 2000 49371
rect 0 49200 2000 49315
rect 0 48765 2000 49000
rect 0 48709 1447 48765
rect 1503 48709 2000 48765
rect 0 48633 2000 48709
rect 0 48577 1447 48633
rect 1503 48577 2000 48633
rect 0 48501 2000 48577
rect 0 48445 1447 48501
rect 1503 48445 2000 48501
rect 0 48369 2000 48445
rect 0 48313 1447 48369
rect 1503 48313 2000 48369
rect 0 48237 2000 48313
rect 0 48181 1447 48237
rect 1503 48181 2000 48237
rect 0 48105 2000 48181
rect 0 48049 1447 48105
rect 1503 48049 2000 48105
rect 0 47973 2000 48049
rect 0 47917 1447 47973
rect 1503 47917 2000 47973
rect 0 47841 2000 47917
rect 0 47785 1447 47841
rect 1503 47785 2000 47841
rect 0 47709 2000 47785
rect 0 47653 1447 47709
rect 1503 47653 2000 47709
rect 0 47577 2000 47653
rect 0 47521 1447 47577
rect 1503 47521 2000 47577
rect 0 47445 2000 47521
rect 0 47389 1447 47445
rect 1503 47389 2000 47445
rect 0 47313 2000 47389
rect 0 47257 1447 47313
rect 1503 47257 2000 47313
rect 0 47181 2000 47257
rect 0 47125 1447 47181
rect 1503 47125 2000 47181
rect 0 47049 2000 47125
rect 0 46993 1447 47049
rect 1503 46993 2000 47049
rect 0 46917 2000 46993
rect 0 46861 1447 46917
rect 1503 46861 2000 46917
rect 0 46785 2000 46861
rect 0 46729 1447 46785
rect 1503 46729 2000 46785
rect 0 46653 2000 46729
rect 0 46597 1447 46653
rect 1503 46597 2000 46653
rect 0 46521 2000 46597
rect 0 46465 1447 46521
rect 1503 46465 2000 46521
rect 0 46389 2000 46465
rect 0 46333 1447 46389
rect 1503 46333 2000 46389
rect 0 46257 2000 46333
rect 0 46201 1447 46257
rect 1503 46201 2000 46257
rect 0 46000 2000 46201
rect 0 45541 2000 45800
rect 0 45485 524 45541
rect 580 45485 2000 45541
rect 0 45409 2000 45485
rect 0 45353 524 45409
rect 580 45353 2000 45409
rect 0 45277 2000 45353
rect 0 45221 524 45277
rect 580 45221 2000 45277
rect 0 45145 2000 45221
rect 0 45089 524 45145
rect 580 45089 2000 45145
rect 0 45013 2000 45089
rect 0 44957 524 45013
rect 580 44957 2000 45013
rect 0 44881 2000 44957
rect 0 44825 524 44881
rect 580 44825 2000 44881
rect 0 44749 2000 44825
rect 0 44693 524 44749
rect 580 44693 2000 44749
rect 0 44617 2000 44693
rect 0 44561 524 44617
rect 580 44561 2000 44617
rect 0 44485 2000 44561
rect 0 44429 524 44485
rect 580 44429 2000 44485
rect 0 44353 2000 44429
rect 0 44297 524 44353
rect 580 44297 2000 44353
rect 0 44221 2000 44297
rect 0 44165 524 44221
rect 580 44165 2000 44221
rect 0 44089 2000 44165
rect 0 44033 524 44089
rect 580 44033 2000 44089
rect 0 43957 2000 44033
rect 0 43901 524 43957
rect 580 43901 2000 43957
rect 0 43825 2000 43901
rect 0 43769 524 43825
rect 580 43769 2000 43825
rect 0 43693 2000 43769
rect 0 43637 524 43693
rect 580 43637 2000 43693
rect 0 43561 2000 43637
rect 0 43505 524 43561
rect 580 43505 2000 43561
rect 0 43429 2000 43505
rect 0 43373 524 43429
rect 580 43373 2000 43429
rect 0 43297 2000 43373
rect 0 43241 524 43297
rect 580 43241 2000 43297
rect 0 43165 2000 43241
rect 0 43109 524 43165
rect 580 43109 2000 43165
rect 0 43033 2000 43109
rect 0 42977 524 43033
rect 580 42977 2000 43033
rect 0 42800 2000 42977
rect 0 42456 2000 42600
rect 0 42400 524 42456
rect 580 42400 2000 42456
rect 0 42324 2000 42400
rect 0 42268 524 42324
rect 580 42268 2000 42324
rect 0 42192 2000 42268
rect 0 42136 524 42192
rect 580 42136 2000 42192
rect 0 42060 2000 42136
rect 0 42004 524 42060
rect 580 42004 2000 42060
rect 0 41928 2000 42004
rect 0 41872 524 41928
rect 580 41872 2000 41928
rect 0 41796 2000 41872
rect 0 41740 524 41796
rect 580 41740 2000 41796
rect 0 41664 2000 41740
rect 0 41608 524 41664
rect 580 41608 2000 41664
rect 0 41532 2000 41608
rect 0 41476 524 41532
rect 580 41476 2000 41532
rect 0 41400 2000 41476
rect 0 41344 524 41400
rect 580 41344 2000 41400
rect 0 41200 2000 41344
rect 0 40884 2000 41000
rect 0 40828 1447 40884
rect 1503 40828 2000 40884
rect 0 40752 2000 40828
rect 0 40696 1447 40752
rect 1503 40696 2000 40752
rect 0 40620 2000 40696
rect 0 40564 1447 40620
rect 1503 40564 2000 40620
rect 0 40488 2000 40564
rect 0 40432 1447 40488
rect 1503 40432 2000 40488
rect 0 40356 2000 40432
rect 0 40300 1447 40356
rect 1503 40300 2000 40356
rect 0 40224 2000 40300
rect 0 40168 1447 40224
rect 1503 40168 2000 40224
rect 0 40092 2000 40168
rect 0 40036 1447 40092
rect 1503 40036 2000 40092
rect 0 39960 2000 40036
rect 0 39904 1447 39960
rect 1503 39904 2000 39960
rect 0 39828 2000 39904
rect 0 39772 1447 39828
rect 1503 39772 2000 39828
rect 0 39600 2000 39772
rect 0 39220 2000 39400
rect 0 39164 524 39220
rect 580 39164 2000 39220
rect 0 39088 2000 39164
rect 0 39032 524 39088
rect 580 39032 2000 39088
rect 0 38956 2000 39032
rect 0 38900 524 38956
rect 580 38900 2000 38956
rect 0 38824 2000 38900
rect 0 38768 524 38824
rect 580 38768 2000 38824
rect 0 38692 2000 38768
rect 0 38636 524 38692
rect 580 38636 2000 38692
rect 0 38560 2000 38636
rect 0 38504 524 38560
rect 580 38504 2000 38560
rect 0 38428 2000 38504
rect 0 38372 524 38428
rect 580 38372 2000 38428
rect 0 38296 2000 38372
rect 0 38240 524 38296
rect 580 38240 2000 38296
rect 0 38164 2000 38240
rect 0 38108 524 38164
rect 580 38108 2000 38164
rect 0 38032 2000 38108
rect 0 37976 524 38032
rect 580 37976 2000 38032
rect 0 37900 2000 37976
rect 0 37844 524 37900
rect 580 37844 2000 37900
rect 0 37768 2000 37844
rect 0 37712 524 37768
rect 580 37712 2000 37768
rect 0 37636 2000 37712
rect 0 37580 524 37636
rect 580 37580 2000 37636
rect 0 37504 2000 37580
rect 0 37448 524 37504
rect 580 37448 2000 37504
rect 0 37372 2000 37448
rect 0 37316 524 37372
rect 580 37316 2000 37372
rect 0 37240 2000 37316
rect 0 37184 524 37240
rect 580 37184 2000 37240
rect 0 37108 2000 37184
rect 0 37052 524 37108
rect 580 37052 2000 37108
rect 0 36976 2000 37052
rect 0 36920 524 36976
rect 580 36920 2000 36976
rect 0 36844 2000 36920
rect 0 36788 524 36844
rect 580 36788 2000 36844
rect 0 36712 2000 36788
rect 0 36656 524 36712
rect 580 36656 2000 36712
rect 0 36400 2000 36656
rect 0 35999 2000 36200
rect 0 35943 524 35999
rect 580 35943 2000 35999
rect 0 35867 2000 35943
rect 0 35811 524 35867
rect 580 35811 2000 35867
rect 0 35735 2000 35811
rect 0 35679 524 35735
rect 580 35679 2000 35735
rect 0 35603 2000 35679
rect 0 35547 524 35603
rect 580 35547 2000 35603
rect 0 35471 2000 35547
rect 0 35415 524 35471
rect 580 35415 2000 35471
rect 0 35339 2000 35415
rect 0 35283 524 35339
rect 580 35283 2000 35339
rect 0 35207 2000 35283
rect 0 35151 524 35207
rect 580 35151 2000 35207
rect 0 35075 2000 35151
rect 0 35019 524 35075
rect 580 35019 2000 35075
rect 0 34943 2000 35019
rect 0 34887 524 34943
rect 580 34887 2000 34943
rect 0 34811 2000 34887
rect 0 34755 524 34811
rect 580 34755 2000 34811
rect 0 34679 2000 34755
rect 0 34623 524 34679
rect 580 34623 2000 34679
rect 0 34547 2000 34623
rect 0 34491 524 34547
rect 580 34491 2000 34547
rect 0 34415 2000 34491
rect 0 34359 524 34415
rect 580 34359 2000 34415
rect 0 34283 2000 34359
rect 0 34227 524 34283
rect 580 34227 2000 34283
rect 0 34151 2000 34227
rect 0 34095 524 34151
rect 580 34095 2000 34151
rect 0 34019 2000 34095
rect 0 33963 524 34019
rect 580 33963 2000 34019
rect 0 33887 2000 33963
rect 0 33831 524 33887
rect 580 33831 2000 33887
rect 0 33755 2000 33831
rect 0 33699 524 33755
rect 580 33699 2000 33755
rect 0 33623 2000 33699
rect 0 33567 524 33623
rect 580 33567 2000 33623
rect 0 33491 2000 33567
rect 0 33435 524 33491
rect 580 33435 2000 33491
rect 0 33200 2000 33435
rect 0 32774 2000 33000
rect 0 32718 524 32774
rect 580 32718 2000 32774
rect 0 32642 2000 32718
rect 0 32586 524 32642
rect 580 32586 2000 32642
rect 0 32510 2000 32586
rect 0 32454 524 32510
rect 580 32454 2000 32510
rect 0 32378 2000 32454
rect 0 32322 524 32378
rect 580 32322 2000 32378
rect 0 32246 2000 32322
rect 0 32190 524 32246
rect 580 32190 2000 32246
rect 0 32114 2000 32190
rect 0 32058 524 32114
rect 580 32058 2000 32114
rect 0 31982 2000 32058
rect 0 31926 524 31982
rect 580 31926 2000 31982
rect 0 31850 2000 31926
rect 0 31794 524 31850
rect 580 31794 2000 31850
rect 0 31718 2000 31794
rect 0 31662 524 31718
rect 580 31662 2000 31718
rect 0 31586 2000 31662
rect 0 31530 524 31586
rect 580 31530 2000 31586
rect 0 31454 2000 31530
rect 0 31398 524 31454
rect 580 31398 2000 31454
rect 0 31322 2000 31398
rect 0 31266 524 31322
rect 580 31266 2000 31322
rect 0 31190 2000 31266
rect 0 31134 524 31190
rect 580 31134 2000 31190
rect 0 31058 2000 31134
rect 0 31002 524 31058
rect 580 31002 2000 31058
rect 0 30926 2000 31002
rect 0 30870 524 30926
rect 580 30870 2000 30926
rect 0 30794 2000 30870
rect 0 30738 524 30794
rect 580 30738 2000 30794
rect 0 30662 2000 30738
rect 0 30606 524 30662
rect 580 30606 2000 30662
rect 0 30530 2000 30606
rect 0 30474 524 30530
rect 580 30474 2000 30530
rect 0 30398 2000 30474
rect 0 30342 524 30398
rect 580 30342 2000 30398
rect 0 30266 2000 30342
rect 0 30210 524 30266
rect 580 30210 2000 30266
rect 0 30000 2000 30210
rect 0 29632 2000 29800
rect 0 29576 524 29632
rect 580 29576 2000 29632
rect 0 29500 2000 29576
rect 0 29444 524 29500
rect 580 29444 2000 29500
rect 0 29368 2000 29444
rect 0 29312 524 29368
rect 580 29312 2000 29368
rect 0 29236 2000 29312
rect 0 29180 524 29236
rect 580 29180 2000 29236
rect 0 29104 2000 29180
rect 0 29048 524 29104
rect 580 29048 2000 29104
rect 0 28972 2000 29048
rect 0 28916 524 28972
rect 580 28916 2000 28972
rect 0 28840 2000 28916
rect 0 28784 524 28840
rect 580 28784 2000 28840
rect 0 28708 2000 28784
rect 0 28652 524 28708
rect 580 28652 2000 28708
rect 0 28576 2000 28652
rect 0 28520 524 28576
rect 580 28520 2000 28576
rect 0 28444 2000 28520
rect 0 28388 524 28444
rect 580 28388 2000 28444
rect 0 28312 2000 28388
rect 0 28256 524 28312
rect 580 28256 2000 28312
rect 0 28180 2000 28256
rect 0 28124 524 28180
rect 580 28124 2000 28180
rect 0 28048 2000 28124
rect 0 27992 524 28048
rect 580 27992 2000 28048
rect 0 27916 2000 27992
rect 0 27860 524 27916
rect 580 27860 2000 27916
rect 0 27784 2000 27860
rect 0 27728 524 27784
rect 580 27728 2000 27784
rect 0 27652 2000 27728
rect 0 27596 524 27652
rect 580 27596 2000 27652
rect 0 27520 2000 27596
rect 0 27464 524 27520
rect 580 27464 2000 27520
rect 0 27388 2000 27464
rect 0 27332 524 27388
rect 580 27332 2000 27388
rect 0 27256 2000 27332
rect 0 27200 524 27256
rect 580 27200 2000 27256
rect 0 27124 2000 27200
rect 0 27068 524 27124
rect 580 27068 2000 27124
rect 0 26800 2000 27068
rect 0 26490 2000 26600
rect 0 26434 1447 26490
rect 1503 26434 2000 26490
rect 0 26358 2000 26434
rect 0 26302 1447 26358
rect 1503 26302 2000 26358
rect 0 26226 2000 26302
rect 0 26170 1447 26226
rect 1503 26170 2000 26226
rect 0 26094 2000 26170
rect 0 26038 1447 26094
rect 1503 26038 2000 26094
rect 0 25962 2000 26038
rect 0 25906 1447 25962
rect 1503 25906 2000 25962
rect 0 25830 2000 25906
rect 0 25774 1447 25830
rect 1503 25774 2000 25830
rect 0 25698 2000 25774
rect 0 25642 1447 25698
rect 1503 25642 2000 25698
rect 0 25566 2000 25642
rect 0 25510 1447 25566
rect 1503 25510 2000 25566
rect 0 25434 2000 25510
rect 0 25378 1447 25434
rect 1503 25378 2000 25434
rect 0 25200 2000 25378
rect 0 24857 2000 25000
rect 0 24801 524 24857
rect 580 24801 2000 24857
rect 0 24725 2000 24801
rect 0 24669 524 24725
rect 580 24669 2000 24725
rect 0 24593 2000 24669
rect 0 24537 524 24593
rect 580 24537 2000 24593
rect 0 24461 2000 24537
rect 0 24405 524 24461
rect 580 24405 2000 24461
rect 0 24329 2000 24405
rect 0 24273 524 24329
rect 580 24273 2000 24329
rect 0 24197 2000 24273
rect 0 24141 524 24197
rect 580 24141 2000 24197
rect 0 24065 2000 24141
rect 0 24009 524 24065
rect 580 24009 2000 24065
rect 0 23933 2000 24009
rect 0 23877 524 23933
rect 580 23877 2000 23933
rect 0 23801 2000 23877
rect 0 23745 524 23801
rect 580 23745 2000 23801
rect 0 23600 2000 23745
rect 0 23151 2000 23400
rect 0 23095 1447 23151
rect 1503 23095 2000 23151
rect 0 23019 2000 23095
rect 0 22963 1447 23019
rect 1503 22963 2000 23019
rect 0 22887 2000 22963
rect 0 22831 1447 22887
rect 1503 22831 2000 22887
rect 0 22755 2000 22831
rect 0 22699 1447 22755
rect 1503 22699 2000 22755
rect 0 22623 2000 22699
rect 0 22567 1447 22623
rect 1503 22567 2000 22623
rect 0 22491 2000 22567
rect 0 22435 1447 22491
rect 1503 22435 2000 22491
rect 0 22359 2000 22435
rect 0 22303 1447 22359
rect 1503 22303 2000 22359
rect 0 22227 2000 22303
rect 0 22171 1447 22227
rect 1503 22171 2000 22227
rect 0 22095 2000 22171
rect 0 22039 1447 22095
rect 1503 22039 2000 22095
rect 0 21963 2000 22039
rect 0 21907 1447 21963
rect 1503 21907 2000 21963
rect 0 21831 2000 21907
rect 0 21775 1447 21831
rect 1503 21775 2000 21831
rect 0 21699 2000 21775
rect 0 21643 1447 21699
rect 1503 21643 2000 21699
rect 0 21567 2000 21643
rect 0 21511 1447 21567
rect 1503 21511 2000 21567
rect 0 21435 2000 21511
rect 0 21379 1447 21435
rect 1503 21379 2000 21435
rect 0 21303 2000 21379
rect 0 21247 1447 21303
rect 1503 21247 2000 21303
rect 0 21171 2000 21247
rect 0 21115 1447 21171
rect 1503 21115 2000 21171
rect 0 21039 2000 21115
rect 0 20983 1447 21039
rect 1503 20983 2000 21039
rect 0 20907 2000 20983
rect 0 20851 1447 20907
rect 1503 20851 2000 20907
rect 0 20775 2000 20851
rect 0 20719 1447 20775
rect 1503 20719 2000 20775
rect 0 20643 2000 20719
rect 0 20587 1447 20643
rect 1503 20587 2000 20643
rect 0 20400 2000 20587
rect 0 20004 2000 20200
rect 0 19948 1447 20004
rect 1503 19948 2000 20004
rect 0 19872 2000 19948
rect 0 19816 1447 19872
rect 1503 19816 2000 19872
rect 0 19740 2000 19816
rect 0 19684 1447 19740
rect 1503 19684 2000 19740
rect 0 19608 2000 19684
rect 0 19552 1447 19608
rect 1503 19552 2000 19608
rect 0 19476 2000 19552
rect 0 19420 1447 19476
rect 1503 19420 2000 19476
rect 0 19344 2000 19420
rect 0 19288 1447 19344
rect 1503 19288 2000 19344
rect 0 19212 2000 19288
rect 0 19156 1447 19212
rect 1503 19156 2000 19212
rect 0 19080 2000 19156
rect 0 19024 1447 19080
rect 1503 19024 2000 19080
rect 0 18948 2000 19024
rect 0 18892 1447 18948
rect 1503 18892 2000 18948
rect 0 18816 2000 18892
rect 0 18760 1447 18816
rect 1503 18760 2000 18816
rect 0 18684 2000 18760
rect 0 18628 1447 18684
rect 1503 18628 2000 18684
rect 0 18552 2000 18628
rect 0 18496 1447 18552
rect 1503 18496 2000 18552
rect 0 18420 2000 18496
rect 0 18364 1447 18420
rect 1503 18364 2000 18420
rect 0 18288 2000 18364
rect 0 18232 1447 18288
rect 1503 18232 2000 18288
rect 0 18156 2000 18232
rect 0 18100 1447 18156
rect 1503 18100 2000 18156
rect 0 18024 2000 18100
rect 0 17968 1447 18024
rect 1503 17968 2000 18024
rect 0 17892 2000 17968
rect 0 17836 1447 17892
rect 1503 17836 2000 17892
rect 0 17760 2000 17836
rect 0 17704 1447 17760
rect 1503 17704 2000 17760
rect 0 17628 2000 17704
rect 0 17572 1447 17628
rect 1503 17572 2000 17628
rect 0 17496 2000 17572
rect 0 17440 1447 17496
rect 1503 17440 2000 17496
rect 0 17200 2000 17440
rect 0 16814 2000 17000
rect 0 16758 1447 16814
rect 1503 16758 2000 16814
rect 0 16682 2000 16758
rect 0 16626 1447 16682
rect 1503 16626 2000 16682
rect 0 16550 2000 16626
rect 0 16494 1447 16550
rect 1503 16494 2000 16550
rect 0 16418 2000 16494
rect 0 16362 1447 16418
rect 1503 16362 2000 16418
rect 0 16286 2000 16362
rect 0 16230 1447 16286
rect 1503 16230 2000 16286
rect 0 16154 2000 16230
rect 0 16098 1447 16154
rect 1503 16098 2000 16154
rect 0 16022 2000 16098
rect 0 15966 1447 16022
rect 1503 15966 2000 16022
rect 0 15890 2000 15966
rect 0 15834 1447 15890
rect 1503 15834 2000 15890
rect 0 15758 2000 15834
rect 0 15702 1447 15758
rect 1503 15702 2000 15758
rect 0 15626 2000 15702
rect 0 15570 1447 15626
rect 1503 15570 2000 15626
rect 0 15494 2000 15570
rect 0 15438 1447 15494
rect 1503 15438 2000 15494
rect 0 15362 2000 15438
rect 0 15306 1447 15362
rect 1503 15306 2000 15362
rect 0 15230 2000 15306
rect 0 15174 1447 15230
rect 1503 15174 2000 15230
rect 0 15098 2000 15174
rect 0 15042 1447 15098
rect 1503 15042 2000 15098
rect 0 14966 2000 15042
rect 0 14910 1447 14966
rect 1503 14910 2000 14966
rect 0 14834 2000 14910
rect 0 14778 1447 14834
rect 1503 14778 2000 14834
rect 0 14702 2000 14778
rect 0 14646 1447 14702
rect 1503 14646 2000 14702
rect 0 14570 2000 14646
rect 0 14514 1447 14570
rect 1503 14514 2000 14570
rect 0 14438 2000 14514
rect 0 14382 1447 14438
rect 1503 14382 2000 14438
rect 0 14306 2000 14382
rect 0 14250 1447 14306
rect 1503 14250 2000 14306
rect 0 14000 2000 14250
use POLY_SUB_FILL_1  POLY_SUB_FILL_1_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
array 0 0 -1950 0 15 3412
timestamp 1765501852
transform -1 0 2287 0 1 14392
box 310 -127 2260 3485
<< labels >>
rlabel metal3 s 1011 50023 1011 50023 4 VSS
port 1 nsew
rlabel metal3 s 1011 64258 1011 64258 4 VSS
port 1 nsew
rlabel metal3 s 1011 62823 1011 62823 4 VDD
port 2 nsew
rlabel metal3 s 1011 51458 1011 51458 4 VDD
port 2 nsew
rlabel metal3 s 1011 69049 1011 69049 4 DVSS
port 3 nsew
rlabel metal3 s 1011 66023 1011 66023 4 DVSS
port 3 nsew
rlabel metal3 s 1011 61058 1011 61058 4 DVSS
port 3 nsew
rlabel metal3 s 1011 57858 1011 57858 4 DVSS
port 3 nsew
rlabel metal3 s 1011 47595 1011 47595 4 DVSS
port 3 nsew
rlabel metal3 s 1011 40342 1011 40342 4 DVSS
port 3 nsew
rlabel metal3 s 1011 26100 1011 26100 4 DVSS
port 3 nsew
rlabel metal3 s 1011 21907 1011 21907 4 DVSS
port 3 nsew
rlabel metal3 s 1011 15750 1011 15750 4 DVSS
port 3 nsew
rlabel metal3 s 1011 18921 1011 18921 4 DVSS
port 3 nsew
rlabel metal3 s 1011 24284 1011 24284 4 DVDD
port 4 nsew
rlabel metal3 s 1011 28394 1011 28394 4 DVDD
port 4 nsew
rlabel metal3 s 1011 31609 1011 31609 4 DVDD
port 4 nsew
rlabel metal3 s 1011 34723 1011 34723 4 DVDD
port 4 nsew
rlabel metal3 s 1011 37959 1011 37959 4 DVDD
port 4 nsew
rlabel metal3 s 1011 41977 1011 41977 4 DVDD
port 4 nsew
rlabel metal3 s 1011 44368 1011 44368 4 DVDD
port 4 nsew
rlabel metal3 s 1011 53223 1011 53223 4 DVDD
port 4 nsew
rlabel metal3 s 1011 54658 1011 54658 4 DVDD
port 4 nsew
rlabel metal3 s 1011 56423 1011 56423 4 DVDD
port 4 nsew
rlabel metal3 s 1011 59623 1011 59623 4 DVDD
port 4 nsew
rlabel metal3 s 1011 67458 1011 67458 4 DVDD
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 2000 70000
<< end >>
