magic
tech gf180mcuD
magscale 1 10
timestamp 1765308861
<< error_p >>
rect -808 -255 -778 -209
rect -594 -255 -564 -209
rect -380 -255 -350 -209
rect -166 -255 -136 -209
rect 53 -255 83 -209
rect 267 -255 297 -209
rect 481 -255 511 -209
rect 695 -255 725 -209
<< nwell >>
rect -1128 -486 1121 486
<< hvpmos >>
rect -810 -176 -700 224
rect -596 -176 -486 224
rect -382 -176 -272 224
rect -168 -176 -58 224
rect 51 -176 161 224
rect 265 -176 375 224
rect 479 -176 589 224
rect 693 -176 803 224
<< mvpdiff >>
rect -898 188 -810 224
rect -898 -140 -885 188
rect -839 -140 -810 188
rect -898 -176 -810 -140
rect -700 188 -596 224
rect -700 -140 -671 188
rect -625 -140 -596 188
rect -700 -176 -596 -140
rect -486 188 -382 224
rect -486 -140 -457 188
rect -411 -140 -382 188
rect -486 -176 -382 -140
rect -272 188 -168 224
rect -272 -140 -243 188
rect -197 -140 -168 188
rect -272 -176 -168 -140
rect -58 188 51 224
rect -58 -140 -29 188
rect 17 -140 51 188
rect -58 -176 51 -140
rect 161 188 265 224
rect 161 -140 190 188
rect 236 -140 265 188
rect 161 -176 265 -140
rect 375 188 479 224
rect 375 -140 404 188
rect 450 -140 479 188
rect 375 -176 479 -140
rect 589 188 693 224
rect 589 -140 618 188
rect 664 -140 693 188
rect 589 -176 693 -140
rect 803 188 891 224
rect 803 -140 832 188
rect 878 -140 891 188
rect 803 -176 891 -140
<< mvpdiffc >>
rect -885 -140 -839 188
rect -671 -140 -625 188
rect -457 -140 -411 188
rect -243 -140 -197 188
rect -29 -140 17 188
rect 190 -140 236 188
rect 404 -140 450 188
rect 618 -140 664 188
rect 832 -140 878 188
<< mvnsubdiff >>
rect -1042 387 1035 400
rect -1042 341 -869 387
rect 869 341 1035 387
rect -1042 328 1035 341
rect -1042 258 -970 328
rect -1042 -258 -1029 258
rect -983 -258 -970 258
rect 963 258 1035 328
rect -1042 -328 -970 -258
rect 963 -258 976 258
rect 1022 -258 1035 258
rect 963 -328 1035 -258
rect -1042 -400 1035 -328
<< mvnsubdiffcont >>
rect -869 341 869 387
rect -1029 -258 -983 258
rect 976 -258 1022 258
<< polysilicon >>
rect -810 224 -700 268
rect -596 224 -486 268
rect -382 224 -272 268
rect -168 224 -58 268
rect 51 224 161 268
rect 265 224 375 268
rect 479 224 589 268
rect 693 224 803 268
rect -810 -209 -700 -176
rect -810 -255 -778 -209
rect -732 -255 -700 -209
rect -810 -268 -700 -255
rect -596 -209 -486 -176
rect -596 -255 -564 -209
rect -518 -255 -486 -209
rect -596 -268 -486 -255
rect -382 -209 -272 -176
rect -382 -255 -350 -209
rect -304 -255 -272 -209
rect -382 -268 -272 -255
rect -168 -209 -58 -176
rect -168 -255 -136 -209
rect -90 -255 -58 -209
rect -168 -268 -58 -255
rect 51 -209 161 -176
rect 51 -255 83 -209
rect 129 -255 161 -209
rect 51 -268 161 -255
rect 265 -209 375 -176
rect 265 -255 297 -209
rect 343 -255 375 -209
rect 265 -268 375 -255
rect 479 -209 589 -176
rect 479 -255 511 -209
rect 557 -255 589 -209
rect 479 -268 589 -255
rect 693 -209 803 -176
rect 693 -255 725 -209
rect 771 -255 803 -209
rect 693 -268 803 -255
<< polycontact >>
rect -778 -255 -732 -209
rect -564 -255 -518 -209
rect -350 -255 -304 -209
rect -136 -255 -90 -209
rect 83 -255 129 -209
rect 297 -255 343 -209
rect 511 -255 557 -209
rect 725 -255 771 -209
<< metal1 >>
rect -1029 341 -869 387
rect 869 341 1022 387
rect -1029 258 -983 341
rect 976 258 1022 341
rect -885 188 -839 222
rect -885 -174 -839 -140
rect -671 188 -625 222
rect -671 -174 -625 -140
rect -457 188 -411 222
rect -457 -174 -411 -140
rect -243 188 -197 222
rect -243 -174 -197 -140
rect -29 188 17 222
rect -29 -174 17 -140
rect 190 188 236 222
rect 190 -174 236 -140
rect 404 188 450 222
rect 404 -174 450 -140
rect 618 188 664 222
rect 618 -174 664 -140
rect 832 188 878 222
rect 832 -174 878 -140
rect -808 -255 -778 -209
rect -732 -255 -702 -209
rect -594 -255 -564 -209
rect -518 -255 -488 -209
rect -380 -255 -350 -209
rect -304 -255 -274 -209
rect -166 -255 -136 -209
rect -90 -255 -60 -209
rect 53 -255 83 -209
rect 129 -255 159 -209
rect 267 -255 297 -209
rect 343 -255 373 -209
rect 481 -255 511 -209
rect 557 -255 587 -209
rect 695 -255 725 -209
rect 771 -255 801 -209
rect -1029 -341 -983 -258
rect 976 -341 1022 -258
rect -1029 -387 1022 -341
<< properties >>
string FIXED_BBOX -960 -364 960 364
string GDS_END 91898
string GDS_FILE ../gds/simple_por.gds.gz
string GDS_START 83958
<< end >>
