magic
tech gf180mcuD
magscale 1 10
timestamp 1765222409
<< metal1 >>
rect -1244 14345 -152 14464
rect 33 14345 4794 14464
rect 4979 14345 7687 14464
rect 7872 14345 8533 14464
rect -1244 14344 8533 14345
rect 9588 13941 9847 14003
rect 11152 13940 11411 14002
rect -1276 13560 -977 13680
rect -854 13560 -380 13680
rect 2459 13561 2474 13680
rect 2659 13561 2676 13680
rect 2459 13560 2676 13561
rect 5899 13561 5921 13680
rect 6106 13561 6129 13680
rect 5899 13560 6129 13561
rect -1276 12776 -380 12896
rect -167 12777 -152 12896
rect 33 12777 50 12896
rect -167 12776 50 12777
rect 4826 12777 4848 12896
rect 5033 12777 5056 12896
rect 4826 12776 5056 12777
rect 7805 12777 7827 12896
rect 8012 12777 8035 12896
rect 7805 12776 8035 12777
rect 2839 11993 2854 12112
rect 3039 11993 3056 12112
rect 2839 11992 3056 11993
rect 5899 11993 5921 12112
rect 6106 11993 6129 12112
rect 5899 11992 6129 11993
rect 11244 11993 11260 12112
rect 11445 11993 11468 12112
rect 11244 11992 11468 11993
rect -167 11209 -152 11328
rect 33 11209 50 11328
rect -167 11208 50 11209
rect 4826 11209 4848 11328
rect 5033 11209 5056 11328
rect 4826 11208 5056 11209
rect 7805 11209 7827 11328
rect 8012 11209 8035 11328
rect 7805 11208 8035 11209
rect 2839 10425 2854 10544
rect 3039 10425 3056 10544
rect 2839 10424 3056 10425
rect 5899 10425 5921 10544
rect 6106 10425 6129 10544
rect 5899 10424 6129 10425
rect 11244 10425 11260 10544
rect 11445 10425 11468 10544
rect 11244 10424 11468 10425
rect -167 9641 -152 9760
rect 33 9641 50 9760
rect -167 9640 50 9641
rect 4826 9641 4848 9760
rect 5033 9641 5056 9760
rect 4826 9640 5056 9641
rect 7805 9641 7827 9760
rect 8012 9641 8035 9760
rect 7805 9640 8035 9641
rect 2839 8857 2854 8976
rect 3039 8857 3056 8976
rect 2839 8856 3056 8857
rect 5899 8857 5921 8976
rect 6106 8857 6129 8976
rect 5899 8856 6129 8857
rect 11244 8857 11260 8976
rect 11445 8857 11468 8976
rect 11244 8856 11468 8857
rect -167 8073 -152 8192
rect 33 8073 50 8192
rect -167 8072 50 8073
rect 4826 8073 4848 8192
rect 5033 8073 5056 8192
rect 4826 8072 5056 8073
rect 7805 8073 7827 8192
rect 8012 8073 8035 8192
rect 7805 8072 8035 8073
rect 2839 7289 2854 7408
rect 3039 7289 3056 7408
rect 2839 7288 3056 7289
rect 5899 7289 5921 7408
rect 6106 7289 6129 7408
rect 5899 7288 6129 7289
rect 11244 7289 11260 7408
rect 11445 7289 11468 7408
rect 11244 7288 11468 7289
rect -167 6505 -152 6624
rect 33 6505 50 6624
rect -167 6504 50 6505
rect 4826 6505 4848 6624
rect 5033 6505 5056 6624
rect 4826 6504 5056 6505
rect 7805 6505 7827 6624
rect 8012 6505 8035 6624
rect 7805 6504 8035 6505
rect 2839 5721 2854 5840
rect 3039 5721 3056 5840
rect 2839 5720 3056 5721
rect 5899 5721 5921 5840
rect 6106 5721 6129 5840
rect 5899 5720 6129 5721
rect 11244 5721 11260 5840
rect 11445 5721 11468 5840
rect 11244 5720 11468 5721
rect -167 4937 -152 5056
rect 33 4937 50 5056
rect -167 4936 50 4937
rect 4826 4937 4848 5056
rect 5033 4937 5056 5056
rect 4826 4936 5056 4937
rect 7805 4937 7827 5056
rect 8012 4937 8035 5056
rect 7805 4936 8035 4937
rect 2839 4153 2854 4272
rect 3039 4153 3056 4272
rect 2839 4152 3056 4153
rect 5899 4153 5921 4272
rect 6106 4153 6129 4272
rect 5899 4152 6129 4153
rect 11225 4153 11260 4272
rect 11445 4153 11486 4272
rect 11225 4152 11486 4153
rect -167 3369 -152 3488
rect 33 3369 50 3488
rect -167 3368 50 3369
rect 4826 3369 4848 3488
rect 5033 3369 5056 3488
rect 4826 3368 5056 3369
rect 7805 3369 7827 3488
rect 8012 3369 8035 3488
rect 7805 3368 8035 3369
<< via1 >>
rect -152 14345 33 14464
rect 4794 14345 4979 14464
rect 7687 14345 7872 14464
rect 8742 13927 8794 14284
rect 9975 13938 10027 14045
rect 10311 13918 10363 14275
rect 11535 13938 11587 14045
rect 11762 13899 11814 14067
rect 2474 13561 2659 13680
rect 5921 13561 6106 13680
rect -152 12777 33 12896
rect 4848 12777 5033 12896
rect 7827 12777 8012 12896
rect 2854 11993 3039 12112
rect 5921 11993 6106 12112
rect 11260 11993 11445 12112
rect -152 11209 33 11328
rect 4848 11209 5033 11328
rect 7827 11209 8012 11328
rect 2854 10425 3039 10544
rect 5921 10425 6106 10544
rect 11260 10425 11445 10544
rect -152 9641 33 9760
rect 4848 9641 5033 9760
rect 7827 9641 8012 9760
rect 2854 8857 3039 8976
rect 5921 8857 6106 8976
rect 11260 8857 11445 8976
rect -152 8073 33 8192
rect 4848 8073 5033 8192
rect 7827 8073 8012 8192
rect 2854 7289 3039 7408
rect 5921 7289 6106 7408
rect 11260 7289 11445 7408
rect -152 6505 33 6624
rect 4848 6505 5033 6624
rect 7827 6505 8012 6624
rect 2854 5721 3039 5840
rect 5921 5721 6106 5840
rect 11260 5721 11445 5840
rect -152 4937 33 5056
rect 4848 4937 5033 5056
rect 7827 4937 8012 5056
rect 2854 4153 3039 4272
rect 5921 4153 6106 4272
rect 11260 4153 11445 4272
rect -152 3369 33 3488
rect 4848 3369 5033 3488
rect 7827 3369 8012 3488
<< metal2 >>
rect -167 14464 50 14466
rect -167 14345 -152 14464
rect 33 14345 50 14464
rect -167 14344 50 14345
rect 4779 14464 4992 14466
rect 4779 14345 4794 14464
rect 4979 14345 4992 14464
rect 4779 14344 4992 14345
rect 7674 14464 7886 14467
rect 7674 14345 7687 14464
rect 7872 14345 7886 14464
rect 7674 14344 7886 14345
rect -158 12896 40 14344
rect 2457 13680 2676 13682
rect 2457 13561 2474 13680
rect 2659 13561 2676 13680
rect 2457 13559 2676 13561
rect 1157 13256 1213 13275
rect -167 12777 -152 12896
rect 33 12777 50 12896
rect -167 12776 50 12777
rect -158 11328 40 12776
rect 863 12473 919 12491
rect -167 11209 -152 11328
rect 33 11209 50 11328
rect -167 11208 50 11209
rect -158 9760 40 11208
rect 863 11016 919 12417
rect 1157 11687 1213 13200
rect 2457 12911 2655 13559
rect 2457 12713 3046 12911
rect 4785 12898 4983 14344
rect 5915 13680 6113 13696
rect 5906 13561 5921 13680
rect 6106 13561 6123 13680
rect 5906 13560 6123 13561
rect 4785 12896 5050 12898
rect 4785 12777 4848 12896
rect 5033 12777 5050 12896
rect 4833 12776 5050 12777
rect 2848 12112 3046 12713
rect 4838 12774 5040 12776
rect 2839 11993 2854 12112
rect 3039 11993 3056 12112
rect 2839 11992 3056 11993
rect 1157 11612 1213 11631
rect 863 10932 919 10960
rect 2848 10544 3046 11992
rect 4838 11328 5036 12774
rect 5915 12112 6113 13560
rect 7681 13031 7879 14344
rect 8740 14284 8796 14549
rect 8740 13927 8742 14284
rect 8794 13927 8796 14284
rect 10309 14275 10365 14541
rect 8740 13911 8796 13927
rect 9973 14045 10029 14060
rect 9973 13938 9975 14045
rect 10027 13938 10029 14045
rect 9973 13815 10029 13938
rect 10309 13918 10311 14275
rect 10363 13918 10365 14275
rect 11759 14067 11817 14084
rect 10309 13903 10365 13918
rect 11533 14045 11589 14060
rect 11533 13938 11535 14045
rect 11587 13938 11589 14045
rect 9640 13759 10029 13815
rect 11533 13781 11589 13938
rect 11759 13899 11762 14067
rect 11814 13899 11817 14067
rect 11759 13788 11817 13899
rect 9640 13256 9696 13759
rect 7681 12896 8017 13031
rect 7681 12833 7827 12896
rect 7812 12777 7827 12833
rect 8012 12777 8029 12896
rect 7812 12776 8029 12777
rect 7819 12774 8019 12776
rect 5906 11993 5921 12112
rect 6106 11993 6123 12112
rect 5906 11992 6123 11993
rect 4833 11209 4848 11328
rect 5033 11209 5050 11328
rect 4833 11208 5050 11209
rect 4838 11206 5040 11208
rect 2839 10425 2854 10544
rect 3039 10425 3056 10544
rect 2839 10424 3056 10425
rect 1200 10008 1256 10045
rect -167 9641 -152 9760
rect 33 9641 50 9760
rect -167 9640 50 9641
rect -158 8192 40 9640
rect 872 9337 928 9355
rect -167 8073 -152 8192
rect 33 8073 50 8192
rect -167 8072 50 8073
rect -158 6624 40 8072
rect 872 7880 928 9281
rect 1200 8551 1256 9952
rect 2848 8976 3046 10424
rect 4838 9760 5036 11206
rect 5915 10544 6113 11992
rect 7819 11328 8017 12774
rect 9640 12584 9696 13200
rect 11305 13725 11589 13781
rect 11671 13730 11817 13788
rect 11305 12877 11361 13725
rect 11671 13368 11729 13730
rect 11671 13287 11729 13312
rect 9640 12507 9696 12528
rect 10986 12821 11361 12877
rect 9951 11576 10007 11591
rect 7812 11209 7827 11328
rect 8012 11209 8029 11328
rect 7812 11208 8029 11209
rect 7819 11206 8019 11208
rect 5906 10425 5921 10544
rect 6106 10425 6123 10544
rect 5906 10424 6123 10425
rect 4833 9641 4848 9760
rect 5033 9641 5050 9760
rect 4833 9640 5050 9641
rect 4838 9638 5040 9640
rect 2839 8857 2854 8976
rect 3039 8857 3056 8976
rect 2839 8856 3056 8857
rect 1200 8466 1256 8495
rect 872 7805 928 7824
rect 2848 7408 3046 8856
rect 4838 8192 5036 9638
rect 5915 8976 6113 10424
rect 7819 9760 8017 11206
rect 9666 10905 9722 10926
rect 7812 9641 7827 9760
rect 8012 9641 8029 9760
rect 7812 9640 8029 9641
rect 7819 9638 8019 9640
rect 5906 8857 5921 8976
rect 6106 8857 6123 8976
rect 5906 8856 6123 8857
rect 4833 8073 4848 8192
rect 5033 8073 5050 8192
rect 4833 8072 5050 8073
rect 4838 8070 5040 8072
rect 2839 7289 2854 7408
rect 3039 7289 3056 7408
rect 2839 7288 3056 7289
rect 1210 6872 1266 6890
rect -167 6505 -152 6624
rect 33 6505 50 6624
rect -167 6504 50 6505
rect -158 5056 40 6504
rect 885 6201 941 6234
rect -167 4937 -152 5056
rect 33 4937 50 5056
rect -167 4936 50 4937
rect -158 3488 40 4936
rect 885 4744 941 6145
rect 1210 5415 1266 6816
rect 2848 5840 3046 7288
rect 4838 6624 5036 8070
rect 5915 7408 6113 8856
rect 7819 8192 8017 9638
rect 9666 9448 9722 10849
rect 9951 10119 10007 11520
rect 9951 10051 10007 10063
rect 9666 9367 9722 9392
rect 9640 8440 9696 8458
rect 7812 8073 7827 8192
rect 8012 8073 8029 8192
rect 7812 8072 8029 8073
rect 7819 8070 8019 8072
rect 5906 7289 5921 7408
rect 6106 7289 6123 7408
rect 5906 7288 6123 7289
rect 4833 6505 4848 6624
rect 5033 6505 5050 6624
rect 4833 6504 5050 6505
rect 4838 6502 5040 6504
rect 2839 5721 2854 5840
rect 3039 5721 3056 5840
rect 2839 5720 3056 5721
rect 1210 5346 1266 5359
rect 885 4644 941 4688
rect 2848 4272 3046 5720
rect 3698 5080 3754 5104
rect 4838 5056 5036 6502
rect 5915 5840 6113 7288
rect 7819 6624 8017 8070
rect 9640 6983 9696 8384
rect 9640 6910 9696 6927
rect 9964 7769 10020 7799
rect 7812 6505 7827 6624
rect 8012 6505 8029 6624
rect 7812 6504 8029 6505
rect 7819 6502 8019 6504
rect 5906 5721 5921 5840
rect 6106 5721 6123 5840
rect 5906 5720 6123 5721
rect 2839 4153 2854 4272
rect 3039 4153 3056 4272
rect 2839 4152 3056 4153
rect -167 3369 -152 3488
rect 33 3369 50 3488
rect -167 3368 50 3369
rect -158 3366 40 3368
rect 2848 3367 3046 4152
rect 3698 3848 3754 5024
rect 4833 4937 4848 5056
rect 5033 4937 5050 5056
rect 4833 4936 5050 4937
rect 3698 3778 3754 3792
rect 4838 4934 5040 4936
rect 4838 3488 5036 4934
rect 5915 4272 6113 5720
rect 7819 5056 8017 6502
rect 9964 6312 10020 7713
rect 9964 6204 10020 6256
rect 9573 5304 9629 5323
rect 7812 4937 7827 5056
rect 8012 4937 8029 5056
rect 7812 4936 8029 4937
rect 9573 4968 9629 5248
rect 7819 4934 8019 4936
rect 5906 4153 5921 4272
rect 6106 4153 6123 4272
rect 5906 4152 6123 4153
rect 4833 3369 4848 3488
rect 5033 3369 5050 3488
rect 4833 3368 5050 3369
rect 5915 3368 6113 4152
rect 7819 3488 8017 4934
rect 9573 4891 9629 4912
rect 9951 4633 10007 4667
rect 9951 3736 10007 4577
rect 10986 4633 11042 12821
rect 10986 4550 11042 4577
rect 11247 12112 11462 12144
rect 11247 11993 11260 12112
rect 11445 11993 11462 12112
rect 11247 10544 11462 11993
rect 11247 10425 11260 10544
rect 11445 10425 11462 10544
rect 11247 8976 11462 10425
rect 11247 8857 11260 8976
rect 11445 8857 11462 8976
rect 11247 7408 11462 8857
rect 11247 7289 11260 7408
rect 11445 7289 11462 7408
rect 11247 5840 11462 7289
rect 11247 5721 11260 5840
rect 11445 5721 11462 5840
rect 9951 3668 10007 3680
rect 11247 4272 11462 5721
rect 11247 4153 11260 4272
rect 11445 4153 11462 4272
rect 7812 3369 7827 3488
rect 8012 3369 8029 3488
rect 7812 3368 8029 3369
rect 11247 3368 11462 4153
rect 4842 3366 5040 3368
rect 7821 3366 8019 3368
<< via2 >>
rect 1157 13200 1213 13256
rect 863 12417 919 12473
rect 1157 11631 1213 11687
rect 863 10960 919 11016
rect 9640 13200 9696 13256
rect 1200 9952 1256 10008
rect 872 9281 928 9337
rect 11671 13312 11729 13368
rect 9640 12528 9696 12584
rect 9951 11520 10007 11576
rect 1200 8495 1256 8551
rect 872 7824 928 7880
rect 9666 10849 9722 10905
rect 1210 6816 1266 6872
rect 885 6145 941 6201
rect 9951 10063 10007 10119
rect 9666 9392 9722 9448
rect 9640 8384 9696 8440
rect 1210 5359 1266 5415
rect 885 4688 941 4744
rect 3698 5024 3754 5080
rect 9640 6927 9696 6983
rect 9964 7713 10020 7769
rect 3698 3792 3754 3848
rect 9964 6256 10020 6312
rect 9573 5248 9629 5304
rect 9573 4912 9629 4968
rect 9951 4577 10007 4633
rect 10986 4577 11042 4633
rect 9951 3680 10007 3736
<< metal3 >>
rect 12086 13536 12141 13592
rect 12085 13424 12143 13480
rect 11651 13312 11671 13368
rect 11729 13312 11755 13368
rect 12083 13312 12145 13368
rect 1128 13200 1157 13256
rect 1213 13200 1247 13256
rect 9607 13200 9640 13256
rect 9696 13200 9728 13256
rect 9605 12528 9640 12584
rect 9696 12528 9726 12584
rect 835 12417 863 12473
rect 919 12417 945 12473
rect 12080 12192 12138 12248
rect 12083 12080 12138 12136
rect 12080 11968 12135 12024
rect 12080 11856 12138 11912
rect 1131 11631 1157 11687
rect 1213 11631 1250 11687
rect 9880 11520 9951 11576
rect 10007 11520 10041 11576
rect 845 10960 863 11016
rect 919 10960 1003 11016
rect 9639 10849 9666 10905
rect 9722 10849 9746 10905
rect 12077 10624 12135 10680
rect 12080 10512 12135 10568
rect 12083 10400 12138 10456
rect 12077 10288 12135 10344
rect 9899 10063 9951 10119
rect 10007 10063 10056 10119
rect 1145 9952 1200 10008
rect 1256 9952 1311 10008
rect 9646 9392 9666 9448
rect 9722 9392 9753 9448
rect 835 9281 872 9337
rect 928 9281 986 9337
rect 12080 9056 12138 9112
rect 12083 8944 12138 9000
rect 12080 8832 12135 8888
rect 12080 8720 12138 8776
rect 1154 8495 1200 8551
rect 1256 8495 1320 8551
rect 9607 8384 9640 8440
rect 9696 8384 9743 8440
rect 847 7824 872 7880
rect 928 7824 999 7880
rect 9939 7713 9964 7769
rect 10020 7713 10058 7769
rect 12077 7488 12135 7544
rect 12080 7376 12135 7432
rect 12083 7264 12138 7320
rect 12077 7152 12135 7208
rect 9601 6927 9640 6983
rect 9696 6927 9737 6983
rect 1198 6816 1210 6872
rect 1266 6816 1302 6872
rect 9883 6256 9964 6312
rect 10020 6256 10044 6312
rect 856 6145 885 6201
rect 941 6145 987 6201
rect 12080 5920 12138 5976
rect 12083 5808 12138 5864
rect 12080 5696 12135 5752
rect 12080 5584 12138 5640
rect 1191 5359 1210 5415
rect 1266 5359 1295 5415
rect 9554 5248 9573 5304
rect 9629 5248 9654 5304
rect 3660 5024 3698 5080
rect 3754 5024 5474 5080
rect 5418 4968 5474 5024
rect 5418 4912 9573 4968
rect 9629 4912 9646 4968
rect 866 4688 885 4744
rect 941 4688 1000 4744
rect 9909 4577 9951 4633
rect 10007 4577 10986 4633
rect 11042 4577 11074 4633
rect 12077 4352 12135 4408
rect 12079 4240 12135 4296
rect 12082 4128 12138 4184
rect 12080 4016 12138 4072
rect 2214 3792 3698 3848
rect 3754 3792 3794 3848
rect 9745 3680 9951 3736
rect 10007 3680 10022 3736
use gf180mcu_as_sc_mcu7t3v3__fillcap_4  gf180mcu_as_sc_mcu7t3v3__fillcap_4_0 $PDKPATH/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532246
transform 1 0 -1052 0 1 13620
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fillcap_8  gf180mcu_as_sc_mcu7t3v3__fillcap_8_0 $PDKPATH/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532312
transform 1 0 7404 0 1 13620
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fillcap_8  gf180mcu_as_sc_mcu7t3v3__fillcap_8_1
timestamp 1751532312
transform 1 0 6508 0 1 13620
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fillcap_8  gf180mcu_as_sc_mcu7t3v3__fillcap_8_2
timestamp 1751532312
transform 1 0 5612 0 1 13620
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fillcap_8  gf180mcu_as_sc_mcu7t3v3__fillcap_8_3
timestamp 1751532312
transform 1 0 4716 0 1 13620
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fillcap_8  gf180mcu_as_sc_mcu7t3v3__fillcap_8_4
timestamp 1751532312
transform 1 0 3596 0 1 13620
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fillcap_8  gf180mcu_as_sc_mcu7t3v3__fillcap_8_5
timestamp 1751532312
transform 1 0 2700 0 1 13620
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fillcap_8  gf180mcu_as_sc_mcu7t3v3__fillcap_8_6
timestamp 1751532312
transform 1 0 1804 0 1 13620
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fillcap_8  gf180mcu_as_sc_mcu7t3v3__fillcap_8_7
timestamp 1751532312
transform 1 0 908 0 1 13620
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fillcap_8  gf180mcu_as_sc_mcu7t3v3__fillcap_8_8
timestamp 1751532312
transform 1 0 -212 0 1 13620
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  gf180mcu_as_sc_mcu7t3v3__diode_2_0 $PDKPATH/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532392
transform -1 0 11884 0 1 13620
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  gf180mcu_as_sc_mcu7t3v3__fill_1_0 $PDKPATH/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532423
transform 1 0 -380 0 1 13620
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  gf180mcu_as_sc_mcu7t3v3__fill_2_0 $PDKPATH/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532440
transform 1 0 -604 0 1 13620
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  gf180mcu_as_sc_mcu7t3v3__tap_2_0 $PDKPATH/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1759751540
transform 1 0 8300 0 1 13620
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  gf180mcu_as_sc_mcu7t3v3__tap_2_1
timestamp 1759751540
transform -1 0 12108 0 1 13620
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  gf180mcu_as_sc_mcu7t3v3__tap_2_2
timestamp 1759751540
transform 1 0 4492 0 1 13620
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  gf180mcu_as_sc_mcu7t3v3__tap_2_3
timestamp 1759751540
transform 1 0 684 0 1 13620
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  gf180mcu_as_sc_mcu7t3v3__tap_2_4
timestamp 1759751540
transform 1 0 -1276 0 1 13620
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  ibufp00 $PDKPATH/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532043
transform -1 0 10092 0 1 13620
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  ibufp01 $PDKPATH/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751896485
transform -1 0 9644 0 1 13620
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  ibufp10
timestamp 1751532043
transform -1 0 11660 0 1 13620
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  ibufp11
timestamp 1751896485
transform -1 0 11212 0 1 13620
box -86 -86 1206 870
use delay_stage  id_1
timestamp 1765222409
transform -1 0 10812 0 -1 4202
box -1438 -96 12174 860
use delay_stage  id_2
timestamp 1765222409
transform 1 0 76 0 1 4222
box -1438 -96 12174 860
use delay_stage  id_3
timestamp 1765222409
transform -1 0 10812 0 -1 5770
box -1438 -96 12174 860
use delay_stage  id_4
timestamp 1765222409
transform -1 0 10812 0 1 5790
box -1438 -96 12174 860
use delay_stage  id_5
timestamp 1765222409
transform 1 0 76 0 -1 7338
box -1438 -96 12174 860
use delay_stage  id_6
timestamp 1765222409
transform 1 0 76 0 1 7358
box -1438 -96 12174 860
use delay_stage  id_7
timestamp 1765222409
transform -1 0 10812 0 -1 8906
box -1438 -96 12174 860
use delay_stage  id_8
timestamp 1765222409
transform -1 0 10812 0 1 8926
box -1438 -96 12174 860
use delay_stage  id_9
timestamp 1765222409
transform 1 0 76 0 -1 10474
box -1438 -96 12174 860
use delay_stage  id_10
timestamp 1765222409
transform 1 0 76 0 1 10494
box -1438 -96 12174 860
use delay_stage  id_11
timestamp 1765222409
transform -1 0 10812 0 -1 12042
box -1438 -96 12174 860
use delay_stage  id_12
timestamp 1765222409
transform -1 0 10812 0 1 12062
box -1438 -96 12174 860
use start_stage  iss
timestamp 1765161918
transform 1 0 -808 0 -1 13630
box -554 -76 13058 880
<< labels >>
flabel metal1 -1276 12776 -380 12896 0 FreeSans 480 0 0 0 vdd
port 0 nsew
flabel metal1 -1276 13560 -977 13680 0 FreeSans 480 0 0 0 vss
port 1 nsew
flabel metal3 12083 13312 12145 13368 0 FreeSans 480 0 0 0 reset
port 2 nsew
flabel metal2 9640 13724 9696 13780 0 FreeSans 480 0 0 0 d0
flabel metal3 12083 12080 12138 12136 0 FreeSans 480 0 0 0 trim[0]
port 3 nsew
flabel metal3 12080 10512 12135 10568 0 FreeSans 480 0 0 0 trim[1]
port 4 nsew
flabel metal3 12083 8944 12138 9000 0 FreeSans 480 0 0 0 trim[2]
port 5 nsew
flabel metal3 12080 7376 12135 7432 0 FreeSans 480 0 0 0 trim[3]
port 6 nsew
flabel metal3 12083 5808 12138 5864 0 FreeSans 480 0 0 0 trim[4]
port 7 nsew
flabel metal3 12086 13536 12141 13592 0 FreeSans 480 0 0 0 trim[12]
port 17 nsew
flabel metal3 12080 5696 12135 5752 0 FreeSans 480 0 0 0 trim[7]
port 10 nsew
flabel metal3 12083 7264 12138 7320 0 FreeSans 480 0 0 0 trim[8]
port 11 nsew
flabel metal3 12080 8832 12135 8888 0 FreeSans 480 0 0 0 trim[9]
port 12 nsew
flabel metal3 12083 10400 12138 10456 0 FreeSans 480 0 0 0 trim[10]
port 13 nsew
flabel metal3 12080 11968 12135 12024 0 FreeSans 480 0 0 0 trim[11]
port 14 nsew
flabel metal3 12079 4240 12135 4296 0 FreeSans 480 0 0 0 trim[5]
port 18 nsew
flabel metal3 12082 4128 12138 4184 0 FreeSans 480 0 0 0 trim[6]
port 19 nsew
flabel metal3 12080 12192 12138 12248 0 FreeSans 480 0 0 0 trim[13]
port 21 nsew
flabel metal3 12085 13424 12143 13480 0 FreeSans 480 0 0 0 trim[25]
port 20 nsew
flabel metal3 12077 10624 12135 10680 0 FreeSans 480 0 0 0 trim[14]
port 22 nsew
flabel metal3 12080 9056 12138 9112 0 FreeSans 480 0 0 0 trim[15]
port 23 nsew
flabel metal3 12077 7488 12135 7544 0 FreeSans 480 0 0 0 trim[16]
port 24 nsew
flabel metal3 12080 5920 12138 5976 0 FreeSans 480 0 0 0 trim[17]
port 25 nsew
flabel metal3 12077 4352 12135 4408 0 FreeSans 480 0 0 0 trim[18]
port 26 nsew
flabel metal3 12080 4016 12138 4072 0 FreeSans 480 0 0 0 trim[19]
port 27 nsew
flabel metal3 12080 5584 12138 5640 0 FreeSans 480 0 0 0 trim[20]
port 28 nsew
flabel metal3 12077 7152 12135 7208 0 FreeSans 480 0 0 0 trim[21]
port 29 nsew
flabel metal3 12080 8720 12138 8776 0 FreeSans 480 0 0 0 trim[22]
port 30 nsew
flabel metal3 12077 10288 12135 10344 0 FreeSans 480 0 0 0 trim[23]
port 31 nsew
flabel metal3 12080 11856 12138 11912 0 FreeSans 480 0 0 0 trim[24]
port 32 nsew
flabel metal2 11305 13659 11361 13715 0 FreeSans 480 0 0 0 d6
flabel metal1 9666 13941 9727 14003 0 FreeSans 480 0 0 0 c0
flabel metal1 11241 13940 11302 14002 0 FreeSans 480 0 0 0 c1
flabel metal2 10309 14467 10365 14541 0 FreeSans 480 90 0 0 clockp[1]
port 33 nsew
flabel metal2 8740 14475 8796 14549 0 FreeSans 480 90 0 0 clockp[0]
port 34 nsew
<< end >>
