magic
tech gf180mcuD
magscale 1 10
timestamp 1765550551
<< metal1 >>
rect 106424 103426 107485 103546
rect 90290 103110 92110 103122
rect 106426 103120 106546 103426
rect 90290 103010 90410 103110
rect 90740 103010 92110 103110
rect 90290 103002 92110 103010
rect 105317 103000 106546 103120
rect 106129 102642 107485 102762
rect 90290 102330 92110 102338
rect 106129 102336 106249 102642
rect 90290 102230 90870 102330
rect 91200 102230 92110 102330
rect 90290 102218 92110 102230
rect 105378 102216 106249 102336
rect 106424 101858 107485 101978
rect 90290 101540 92110 101554
rect 106426 101552 106546 101858
rect 90290 101440 90410 101540
rect 90740 101440 92110 101540
rect 90290 101434 92110 101440
rect 105378 101432 106546 101552
rect 106129 101074 107485 101194
rect 90290 100760 92110 100770
rect 106129 100768 106249 101074
rect 90290 100660 90870 100760
rect 91200 100660 92110 100760
rect 90290 100650 92110 100660
rect 105378 100648 106249 100768
rect 106424 100290 107485 100410
rect 90290 99980 92110 99986
rect 106426 99984 106546 100290
rect 90290 99880 90410 99980
rect 90740 99880 92110 99980
rect 90290 99866 92110 99880
rect 105378 99864 106546 99984
rect 106129 99506 107485 99626
rect 90290 99190 92110 99202
rect 106129 99200 106249 99506
rect 90290 99090 90870 99190
rect 91200 99090 92110 99190
rect 90290 99082 92110 99090
rect 105378 99080 106249 99200
rect 106424 98722 107485 98842
rect 90290 98410 92110 98418
rect 106426 98416 106546 98722
rect 90290 98310 90410 98410
rect 90740 98310 92110 98410
rect 90290 98298 92110 98310
rect 105378 98296 106546 98416
rect 106129 97938 107485 98058
rect 90290 97630 92110 97634
rect 106129 97632 106249 97938
rect 90290 97530 90870 97630
rect 91200 97530 92110 97630
rect 90290 97514 92110 97530
rect 105378 97512 106249 97632
rect 106424 97154 107485 97274
rect 90290 96840 92110 96850
rect 106426 96848 106546 97154
rect 90290 96740 90410 96840
rect 90740 96740 92110 96840
rect 90290 96730 92110 96740
rect 105378 96728 106546 96848
rect 106129 96370 107485 96490
rect 90290 96050 92110 96066
rect 106129 96064 106249 96370
rect 90290 95950 90870 96050
rect 91200 95950 92110 96050
rect 90290 95946 92110 95950
rect 105378 95944 106249 96064
rect 106424 95586 107485 95706
rect 90290 95270 92110 95282
rect 106426 95280 106546 95586
rect 90290 95170 90410 95270
rect 90740 95170 92110 95270
rect 90290 95162 92110 95170
rect 105378 95160 106546 95280
rect 106129 94802 107485 94922
rect 90290 94490 92110 94498
rect 106129 94496 106249 94802
rect 90290 94390 90870 94490
rect 91200 94390 92110 94490
rect 90290 94378 92110 94390
rect 105378 94376 106249 94496
rect 106424 94018 107485 94138
rect 90290 93700 92110 93714
rect 106426 93712 106546 94018
rect 90290 93600 90410 93700
rect 90740 93600 92110 93700
rect 90290 93594 92110 93600
rect 105378 93592 106546 93712
rect 106129 93234 107485 93354
rect 90290 92920 92110 92930
rect 106129 92928 106249 93234
rect 90290 92820 90870 92920
rect 91200 92820 92110 92920
rect 90290 92810 92110 92820
rect 105378 92808 106249 92928
rect 106424 92450 107485 92570
rect 90290 92140 92110 92146
rect 106426 92144 106546 92450
rect 90290 92040 90410 92140
rect 90740 92040 92110 92140
rect 90290 92026 92110 92040
rect 105379 92024 106546 92144
<< via1 >>
rect 90410 103010 90740 103110
rect 90870 102230 91200 102330
rect 90410 101440 90740 101540
rect 90870 100660 91200 100760
rect 90410 99880 90740 99980
rect 90870 99090 91200 99190
rect 90410 98310 90740 98410
rect 90870 97530 91200 97630
rect 90410 96740 90740 96840
rect 90870 95950 91200 96050
rect 90410 95170 90740 95270
rect 90870 94390 91200 94490
rect 90410 93600 90740 93700
rect 90870 92820 91200 92920
rect 90410 92040 90740 92140
<< metal2 >>
rect 90400 103110 90750 103220
rect 90400 103010 90410 103110
rect 90740 103010 90750 103110
rect 90400 101979 90750 103010
rect 90400 101540 90750 101859
rect 90400 101440 90410 101540
rect 90740 101440 90750 101540
rect 90400 100411 90750 101440
rect 90400 99980 90750 100291
rect 90400 99880 90410 99980
rect 90740 99880 90750 99980
rect 90400 98843 90750 99880
rect 90400 98410 90750 98723
rect 90400 98310 90410 98410
rect 90740 98310 90750 98410
rect 90400 97275 90750 98310
rect 90400 96840 90750 97155
rect 90400 96740 90410 96840
rect 90740 96740 90750 96840
rect 90400 95707 90750 96740
rect 90400 95270 90750 95587
rect 90400 95170 90410 95270
rect 90740 95170 90750 95270
rect 90400 94139 90750 95170
rect 90400 93700 90750 94019
rect 90400 93600 90410 93700
rect 90740 93600 90750 93700
rect 90400 92571 90750 93600
rect 90400 92140 90750 92451
rect 90400 92040 90410 92140
rect 90740 92040 90750 92140
rect 90400 91940 90750 92040
rect 90860 102775 91210 103220
rect 90860 102330 91210 102635
rect 90860 102230 90870 102330
rect 91200 102230 91210 102330
rect 90860 101207 91210 102230
rect 90860 100760 91210 101067
rect 90860 100660 90870 100760
rect 91200 100660 91210 100760
rect 90860 99639 91210 100660
rect 90860 99190 91210 99499
rect 90860 99090 90870 99190
rect 91200 99090 91210 99190
rect 90860 98071 91210 99090
rect 90860 97630 91210 97931
rect 90860 97530 90870 97630
rect 91200 97530 91210 97630
rect 90860 96503 91210 97530
rect 90860 96050 91210 96363
rect 90860 95950 90870 96050
rect 91200 95950 91210 96050
rect 90860 94935 91210 95950
rect 90860 94490 91210 94795
rect 90860 94390 90870 94490
rect 91200 94390 91210 94490
rect 90860 93367 91210 94390
rect 90860 92920 91210 93227
rect 90860 92820 90870 92920
rect 91200 92820 91210 92920
rect 90860 91940 91210 92820
<< via2 >>
rect 90400 101859 90750 101979
rect 90400 100291 90750 100411
rect 90400 98723 90750 98843
rect 90400 97155 90750 97275
rect 90400 95587 90750 95707
rect 90400 94019 90750 94139
rect 90400 92451 90750 92571
rect 90860 102635 91210 102775
rect 90860 101067 91210 101207
rect 90860 99499 91210 99639
rect 90860 97931 91210 98071
rect 90860 96363 91210 96503
rect 90860 94795 91210 94935
rect 90860 93227 91210 93367
<< metal3 >>
rect 88496 102635 90860 102775
rect 91210 102635 91240 102775
rect 88496 101859 90400 101979
rect 90750 101859 90770 101979
rect 88496 101067 90860 101207
rect 91210 101067 91240 101207
rect 88382 100291 90400 100411
rect 90750 100291 90770 100411
rect 88496 99499 90860 99639
rect 91210 99499 91240 99639
rect 88367 98723 90400 98843
rect 90750 98723 90770 98843
rect 88496 97931 90860 98071
rect 91210 97931 91240 98071
rect 88381 97155 90400 97275
rect 90750 97155 90770 97275
rect 88496 96363 90860 96503
rect 91210 96363 91240 96503
rect 88374 95587 90400 95707
rect 90750 95587 90770 95707
rect 88496 94795 90860 94935
rect 91210 94795 91240 94935
rect 88402 94019 90400 94139
rect 90750 94019 90770 94139
rect 88496 93227 90860 93367
rect 91210 93227 91240 93367
rect 88388 92451 90400 92571
rect 90750 92451 90770 92571
<< end >>
