magic
tech gf180mcuD
magscale 1 10
timestamp 1765308861
<< nwell >>
rect 1353 -110 1490 561
rect 1353 -418 2231 -110
rect 1353 -1211 1490 -418
<< metal1 >>
rect 526 385 3034 685
rect 744 -884 883 385
rect 1072 260 1124 300
rect 1072 -872 1124 -832
rect 946 -996 969 -944
rect 1021 -996 1044 -944
rect 946 -1019 1044 -996
rect 1242 -1112 1614 385
rect 1727 309 1779 310
rect 1706 286 1779 309
rect 1706 234 1727 286
rect 1706 209 1779 234
rect 2237 286 2310 310
rect 2289 234 2310 286
rect 2237 210 2310 234
rect 2400 208 2706 385
rect 1841 165 2166 167
rect 1841 113 1873 165
rect 2133 113 2166 165
rect 1841 111 2166 113
rect 2400 52 2634 208
rect 2686 52 2706 208
rect 2400 -2 2706 52
rect 2808 -62 3008 6
rect 2364 -126 3008 -62
rect 2364 -178 2383 -126
rect 2539 -178 3008 -126
rect 2364 -194 3008 -178
rect 2364 -243 2561 -194
rect 1869 -329 2420 -317
rect 1869 -340 2421 -329
rect 1869 -392 1892 -340
rect 2048 -392 2421 -340
rect 1869 -414 2421 -392
rect 1722 -702 1774 -681
rect 1722 -879 1774 -858
rect 1942 -702 1994 -681
rect 1942 -879 1994 -858
rect 1813 -998 1837 -946
rect 1889 -998 1913 -946
rect 1813 -999 1913 -998
rect 589 -1190 789 -1168
rect 589 -1346 610 -1190
rect 766 -1346 789 -1190
rect 2284 -1304 2421 -414
rect 2595 -429 2767 -425
rect 2595 -481 2653 -429
rect 2705 -481 2767 -429
rect 2595 -484 2767 -481
rect 589 -1568 789 -1346
rect 1072 -1490 1118 -1438
rect 1170 -1490 1214 -1438
rect 877 -2015 1021 -1541
rect 1243 -1613 1297 -1559
rect 1295 -1873 1297 -1613
rect 1243 -1927 1297 -1873
rect 1401 -2015 1625 -1320
rect 1825 -1474 1868 -1422
rect 1920 -1474 1963 -1422
rect 1743 -1548 1795 -1531
rect 1993 -1560 2045 -1531
rect 1993 -1850 2045 -1820
rect 1743 -1930 1795 -1912
rect 2171 -2015 2421 -1304
rect 2514 -597 2566 -568
rect 2514 -1926 2566 -1897
rect 2824 -577 2876 -528
rect 2824 -1926 2876 -1877
rect 607 -2315 3034 -2015
<< via1 >>
rect 1072 -832 1124 260
rect 969 -996 1021 -944
rect 1727 234 1779 286
rect 2237 234 2289 286
rect 1873 113 2133 165
rect 2634 52 2686 208
rect 2383 -178 2539 -126
rect 1892 -392 2048 -340
rect 1722 -858 1774 -702
rect 1942 -858 1994 -702
rect 1837 -998 1889 -946
rect 610 -1346 766 -1190
rect 2653 -481 2705 -429
rect 1118 -1490 1170 -1438
rect 1243 -1873 1295 -1613
rect 1868 -1474 1920 -1422
rect 1743 -1912 1795 -1548
rect 1993 -1820 2045 -1560
rect 2514 -1897 2566 -597
rect 2824 -1877 2876 -577
<< metal2 >>
rect 2242 313 2359 333
rect 1070 303 1126 304
rect 1725 303 1781 313
rect 1070 286 1781 303
rect 1070 260 1727 286
rect 1070 -832 1072 260
rect 1124 234 1727 260
rect 1779 234 1781 286
rect 1124 224 1781 234
rect 1124 -707 1126 224
rect 1725 207 1781 224
rect 2235 286 2359 313
rect 2235 234 2237 286
rect 2289 234 2359 286
rect 2235 207 2359 234
rect 2242 190 2359 207
rect 2622 208 2698 236
rect 1841 165 2166 170
rect 1841 113 1873 165
rect 2133 113 2166 165
rect 1841 109 2166 113
rect 1847 -175 1921 109
rect 2242 52 2318 190
rect 1719 -249 1921 -175
rect 1992 -24 2318 52
rect 2622 52 2634 208
rect 2686 52 2698 208
rect 2622 33 2698 52
rect 1719 -465 1793 -249
rect 1992 -322 2068 -24
rect 2364 -97 2561 -62
rect 2128 -126 2561 -97
rect 2128 -178 2383 -126
rect 2539 -178 2561 -126
rect 2128 -226 2561 -178
rect 1869 -340 2070 -322
rect 1869 -392 1892 -340
rect 2048 -392 2070 -340
rect 1869 -408 2070 -392
rect 2128 -422 2257 -226
rect 2364 -243 2561 -226
rect 2622 -239 2696 33
rect 2622 -317 2889 -239
rect 2128 -429 2764 -422
rect 2128 -465 2653 -429
rect 1719 -481 2653 -465
rect 2705 -481 2764 -429
rect 1719 -486 2764 -481
rect 1719 -539 2257 -486
rect 1720 -702 1776 -680
rect 1720 -707 1722 -702
rect 1124 -832 1722 -707
rect 1070 -855 1722 -832
rect 1070 -876 1126 -855
rect 1720 -858 1722 -855
rect 1774 -858 1776 -702
rect 1720 -880 1776 -858
rect 1940 -687 1996 -680
rect 2128 -687 2257 -539
rect 1940 -702 2257 -687
rect 1940 -858 1942 -702
rect 1994 -853 2257 -702
rect 1994 -858 1996 -853
rect 1940 -880 1996 -858
rect 946 -944 1044 -942
rect 946 -996 969 -944
rect 1021 -996 1044 -944
rect 946 -998 1044 -996
rect 1813 -946 1913 -944
rect 1813 -998 1837 -946
rect 1889 -998 1913 -946
rect 589 -1190 789 -1168
rect 589 -1346 610 -1190
rect 766 -1236 789 -1190
rect 961 -1236 1026 -998
rect 1813 -1000 1913 -998
rect 1832 -1236 1907 -1000
rect 766 -1305 1907 -1236
rect 766 -1346 789 -1305
rect 589 -1368 789 -1346
rect 961 -1421 1026 -1305
rect 1832 -1420 1907 -1305
rect 961 -1438 1215 -1421
rect 961 -1486 1118 -1438
rect 1072 -1490 1118 -1486
rect 1170 -1486 1215 -1438
rect 1825 -1422 1963 -1420
rect 1825 -1474 1868 -1422
rect 1920 -1474 1963 -1422
rect 1825 -1476 1963 -1474
rect 1170 -1490 1214 -1486
rect 1072 -1492 1214 -1490
rect 1741 -1548 1797 -1527
rect 1241 -1613 1297 -1555
rect 1241 -1873 1243 -1613
rect 1295 -1634 1297 -1613
rect 1741 -1634 1743 -1548
rect 1295 -1846 1743 -1634
rect 1295 -1873 1297 -1846
rect 1241 -1931 1297 -1873
rect 1741 -1912 1743 -1846
rect 1795 -1912 1797 -1548
rect 1991 -1557 2047 -1527
rect 2128 -1557 2257 -853
rect 1991 -1560 2257 -1557
rect 1991 -1820 1993 -1560
rect 2045 -1805 2257 -1560
rect 2512 -597 2568 -564
rect 2045 -1820 2047 -1805
rect 1991 -1853 2047 -1820
rect 2512 -1897 2514 -597
rect 2566 -1897 2568 -597
rect 2512 -1912 2568 -1897
rect 1741 -1985 2568 -1912
rect 2822 -577 2889 -317
rect 2822 -1877 2824 -577
rect 2876 -1877 2889 -577
rect 2822 -1926 2889 -1877
rect 2822 -1930 2878 -1926
use nmos_6p0_BJPB5U  nmos_6p0_BJPB5U_0
timestamp 1765308861
transform 1 0 1894 0 1 -1706
box -334 -432 334 432
use pmos_6p0_UXEQNM  pmos_6p0_UXEQNM_0
timestamp 1765308861
transform 1 0 1863 0 1 -804
box -378 -386 368 386
use nmos_6p0_L3YBEV  X6
timestamp 1765308861
transform 1 0 2695 0 1 -1203
box -364 -932 364 932
use pmos_6p0_9YEQN4  XM1
timestamp 1765308861
transform 1 0 985 0 1 -325
box -378 -886 368 886
use nmos_6p0_BJPB5U  XM3
timestamp 1765308861
transform 1 0 1144 0 1 -1704
box -334 -432 334 432
use pmos_6p0_9859UL  XM5
timestamp 1765308861
transform 1 0 2008 0 1 226
box -518 -336 518 336
<< labels >>
flabel metal1 s 577 445 777 645 0 FreeSans 1600 0 0 0 VDD
port 1 nsew
flabel metal1 s 639 -2288 839 -2088 0 FreeSans 1600 0 0 0 VSS
port 2 nsew
flabel metal1 s 589 -1568 789 -1368 0 FreeSans 1600 0 0 0 Vin
port 3 nsew
flabel metal1 s 2808 -194 3008 6 0 FreeSans 1600 0 0 0 Vout
port 4 nsew
<< properties >>
string GDS_END 56978
string GDS_FILE ../gds/simple_por.gds.gz
string GDS_START 45324
<< end >>
