magic
tech gf180mcuD
magscale 1 10
timestamp 1765308861
<< pwell >>
rect -1066 -432 1066 432
<< hvnmos >>
rect -802 -224 -662 176
rect -558 -224 -418 176
rect -314 -224 -174 176
rect -70 -224 70 176
rect 174 -224 314 176
rect 418 -224 558 176
rect 662 -224 802 176
<< mvndiff >>
rect -890 140 -802 176
rect -890 -188 -877 140
rect -831 -188 -802 140
rect -890 -224 -802 -188
rect -662 140 -558 176
rect -662 -188 -633 140
rect -587 -188 -558 140
rect -662 -224 -558 -188
rect -418 140 -314 176
rect -418 -188 -389 140
rect -343 -188 -314 140
rect -418 -224 -314 -188
rect -174 140 -70 176
rect -174 -188 -145 140
rect -99 -188 -70 140
rect -174 -224 -70 -188
rect 70 140 174 176
rect 70 -188 99 140
rect 145 -188 174 140
rect 70 -224 174 -188
rect 314 140 418 176
rect 314 -188 343 140
rect 389 -188 418 140
rect 314 -224 418 -188
rect 558 140 662 176
rect 558 -188 587 140
rect 633 -188 662 140
rect 558 -224 662 -188
rect 802 140 890 176
rect 802 -188 831 140
rect 877 -188 890 140
rect 802 -224 890 -188
<< mvndiffc >>
rect -877 -188 -831 140
rect -633 -188 -587 140
rect -389 -188 -343 140
rect -145 -188 -99 140
rect 99 -188 145 140
rect 343 -188 389 140
rect 587 -188 633 140
rect 831 -188 877 140
<< mvpsubdiff >>
rect -1034 328 1034 400
rect -1034 258 -962 328
rect -1034 -258 -1021 258
rect -975 -258 -962 258
rect 962 258 1034 328
rect -1034 -328 -962 -258
rect 962 -258 975 258
rect 1021 -258 1034 258
rect 962 -328 1034 -258
rect -1034 -341 1034 -328
rect -1034 -387 -916 -341
rect 916 -387 1034 -341
rect -1034 -400 1034 -387
<< mvpsubdiffcont >>
rect -1021 -258 -975 258
rect 975 -258 1021 258
rect -916 -387 916 -341
<< polysilicon >>
rect -802 255 -662 268
rect -802 209 -755 255
rect -709 209 -662 255
rect -802 176 -662 209
rect -558 255 -418 268
rect -558 209 -511 255
rect -465 209 -418 255
rect -558 176 -418 209
rect -314 255 -174 268
rect -314 209 -267 255
rect -221 209 -174 255
rect -314 176 -174 209
rect -70 255 70 268
rect -70 209 -23 255
rect 23 209 70 255
rect -70 176 70 209
rect 174 255 314 268
rect 174 209 221 255
rect 267 209 314 255
rect 174 176 314 209
rect 418 255 558 268
rect 418 209 465 255
rect 511 209 558 255
rect 418 176 558 209
rect 662 255 802 268
rect 662 209 709 255
rect 755 209 802 255
rect 662 176 802 209
rect -802 -268 -662 -224
rect -558 -268 -418 -224
rect -314 -268 -174 -224
rect -70 -268 70 -224
rect 174 -268 314 -224
rect 418 -268 558 -224
rect 662 -268 802 -224
<< polycontact >>
rect -755 209 -709 255
rect -511 209 -465 255
rect -267 209 -221 255
rect -23 209 23 255
rect 221 209 267 255
rect 465 209 511 255
rect 709 209 755 255
<< metal1 >>
rect -1021 341 1021 387
rect -1021 258 -975 341
rect 975 258 1021 341
rect -800 209 -755 255
rect -709 209 -664 255
rect -556 209 -511 255
rect -465 209 -420 255
rect -312 209 -267 255
rect -221 209 -176 255
rect -68 209 -23 255
rect 23 209 68 255
rect 176 209 221 255
rect 267 209 312 255
rect 420 209 465 255
rect 511 209 556 255
rect 664 209 709 255
rect 755 209 800 255
rect -877 140 -831 174
rect -877 -222 -831 -188
rect -633 140 -587 174
rect -633 -222 -587 -188
rect -389 140 -343 174
rect -389 -222 -343 -188
rect -145 140 -99 174
rect -145 -222 -99 -188
rect 99 140 145 174
rect 99 -222 145 -188
rect 343 140 389 174
rect 343 -222 389 -188
rect 587 140 633 174
rect 587 -222 633 -188
rect 831 140 877 174
rect 831 -222 877 -188
rect -1021 -341 -975 -258
rect 975 -341 1021 -258
rect -1021 -387 -916 -341
rect 916 -387 1021 -341
<< properties >>
string FIXED_BBOX -998 -364 998 364
string GDS_END 76412
string GDS_FILE ../gds/simple_por.gds.gz
string GDS_START 68920
<< end >>
