magic
tech gf180mcuD
magscale 1 10
timestamp 1765222409
<< nwell >>
rect 460 344 722 860
<< pwell >>
rect 460 260 722 344
<< metal1 >>
rect -1128 714 -605 834
rect 1639 311 1943 361
rect 4338 416 4340 468
rect 1639 304 1951 311
rect -1128 -70 -605 50
<< via1 >>
rect -1026 261 -974 430
rect 46 308 102 415
rect 200 308 256 415
rect 494 308 550 415
rect 648 308 704 415
rect 942 314 998 421
rect 1943 311 1999 418
rect 2592 314 2648 421
rect 3079 406 3276 458
rect 4340 416 4535 468
rect 5088 409 5285 461
rect 6357 414 6552 466
rect 4218 200 4270 369
rect 6235 200 6287 369
rect 6766 313 6819 411
rect 6921 262 6974 428
rect 7340 407 7537 459
rect 8473 269 8526 435
rect 8597 415 8791 467
rect 9132 403 9329 455
rect 10265 279 10318 445
rect 10391 413 10584 465
rect 11741 250 11794 416
<< metal2 >>
rect 632 690 648 746
rect 704 690 722 746
rect 5110 690 5125 746
rect 5181 690 5199 746
rect -1029 430 -971 445
rect -1029 261 -1026 430
rect -974 261 -971 430
rect 46 425 102 434
rect 200 425 256 436
rect 44 415 104 425
rect 44 308 46 415
rect 102 308 104 415
rect 44 295 104 308
rect 198 415 258 425
rect 198 308 200 415
rect 256 308 258 415
rect 198 298 258 308
rect 198 295 200 298
rect -1029 74 -971 261
rect 46 74 102 295
rect 256 295 258 298
rect 492 415 552 428
rect 648 425 704 690
rect 2592 634 2648 686
rect 942 522 998 534
rect 942 431 998 466
rect 1940 522 2002 535
rect 492 308 494 415
rect 550 308 552 415
rect 492 295 552 308
rect 646 415 706 425
rect 646 308 648 415
rect 704 308 706 415
rect 646 295 706 308
rect 940 421 1000 431
rect 940 314 942 421
rect 998 314 1000 421
rect 940 301 1000 314
rect 1940 418 2002 466
rect 2592 431 2648 578
rect 3129 462 3185 478
rect 3067 458 3289 462
rect 1940 311 1943 418
rect 1999 311 2002 418
rect 200 199 256 242
rect 494 186 550 295
rect 1940 280 2002 311
rect 2590 421 2650 431
rect 2590 314 2592 421
rect 2648 314 2650 421
rect 3067 406 3079 458
rect 3276 406 3289 458
rect 3067 402 3289 406
rect 4216 410 4272 685
rect 4369 634 4425 648
rect 4369 472 4425 578
rect 4328 468 4547 472
rect 4328 416 4340 468
rect 4535 416 4547 468
rect 5125 464 5181 690
rect 10425 634 10481 648
rect 6371 522 6428 560
rect 6345 466 6371 469
rect 6919 522 6976 557
rect 6428 466 6564 469
rect 4328 412 4547 416
rect 5075 461 5303 464
rect 2590 301 2650 314
rect 494 85 550 130
rect 3129 186 3185 402
rect 5075 409 5088 461
rect 5285 409 5303 461
rect 5075 406 5303 409
rect 6232 410 6289 421
rect 6345 414 6357 466
rect 6552 414 6564 466
rect 6345 411 6564 414
rect 6764 411 6821 507
rect 4216 200 4218 354
rect 4270 200 4272 354
rect 4216 188 4272 200
rect 6232 200 6235 354
rect 6287 200 6289 354
rect 6764 410 6766 411
rect 6819 410 6821 411
rect 6764 313 6766 354
rect 6819 313 6821 354
rect 6764 233 6821 313
rect 8724 522 8780 536
rect 6919 428 6976 466
rect 7443 462 7499 476
rect 8585 467 8724 470
rect 8780 467 8806 470
rect 10425 468 10481 578
rect 6919 262 6921 428
rect 6974 262 6976 428
rect 7325 459 7552 462
rect 7325 407 7340 459
rect 7537 407 7552 459
rect 8471 451 8527 457
rect 7325 405 7552 407
rect 8470 435 8529 451
rect 8470 410 8473 435
rect 8526 410 8529 435
rect 8585 415 8597 467
rect 8791 415 8806 467
rect 9175 458 9231 466
rect 10379 465 10596 468
rect 8585 412 8806 415
rect 9119 455 9341 458
rect 6919 250 6976 262
rect 6232 187 6289 200
rect 3129 85 3185 130
rect 7443 74 7499 405
rect 8724 401 8780 412
rect 9119 403 9132 455
rect 9329 403 9341 455
rect 9119 401 9341 403
rect 10262 445 10321 462
rect 10262 410 10265 445
rect 10318 410 10321 445
rect 10379 413 10391 465
rect 10584 413 10596 465
rect 10379 411 10596 413
rect 11738 416 11797 435
rect 8470 269 8473 354
rect 8526 269 8529 354
rect 8470 257 8529 269
rect 9175 298 9231 401
rect 10425 384 10481 411
rect 10262 279 10265 354
rect 10318 279 10321 354
rect 10262 266 10321 279
rect 9175 183 9231 242
rect 11738 250 11741 416
rect 11794 250 11797 416
rect 11738 186 11797 250
rect 11738 117 11797 130
rect -1049 18 -1029 74
rect -971 18 -953 74
rect 33 18 46 74
rect 102 18 114 74
rect 7431 18 7443 74
rect 7499 18 7510 74
<< via2 >>
rect 648 690 704 746
rect 5125 690 5181 746
rect 200 242 256 298
rect 2592 578 2648 634
rect 942 466 998 522
rect 1940 466 2002 522
rect 4369 578 4425 634
rect 10425 578 10481 634
rect 6371 466 6428 522
rect 494 130 550 186
rect 4216 369 4272 410
rect 4216 354 4218 369
rect 4218 354 4270 369
rect 4270 354 4272 369
rect 6232 369 6289 410
rect 6232 354 6235 369
rect 6235 354 6287 369
rect 6287 354 6289 369
rect 6764 354 6766 410
rect 6766 354 6819 410
rect 6819 354 6821 410
rect 6919 466 6976 522
rect 8724 467 8780 522
rect 8724 466 8780 467
rect 3129 130 3185 186
rect 8470 354 8473 410
rect 8473 354 8526 410
rect 8526 354 8529 410
rect 9175 242 9231 298
rect 10262 354 10265 410
rect 10265 354 10318 410
rect 10318 354 10321 410
rect 11738 130 11797 186
rect -1029 18 -971 74
rect 46 18 102 74
rect 7443 18 7499 74
<< metal3 >>
rect 623 690 648 746
rect 704 690 5125 746
rect 5181 690 5199 746
rect 2568 578 2592 634
rect 2648 578 4369 634
rect 4425 578 4437 634
rect 6671 578 10425 634
rect 10481 578 10498 634
rect 6671 522 6727 578
rect 922 466 942 522
rect 998 466 1207 522
rect 1928 466 1940 522
rect 2002 466 6371 522
rect 6428 466 6727 522
rect 6895 466 6919 522
rect 6976 466 8724 522
rect 8780 466 8833 522
rect 4200 354 4216 410
rect 4272 354 6232 410
rect 6289 354 6764 410
rect 6821 354 6866 410
rect 8441 354 8470 410
rect 8529 354 10262 410
rect 10321 354 10334 410
rect 181 242 200 298
rect 256 242 9175 298
rect 9231 242 9258 298
rect -1326 130 494 186
rect 550 130 3129 186
rect 3185 130 11738 186
rect 11797 130 12059 186
rect -1326 18 -1029 74
rect -971 18 46 74
rect 102 18 7443 74
rect 7499 18 12059 74
use gf180mcu_as_sc_mcu7t3v3__invz_2  delanenb0 $PDKPATH/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1764933398
transform 1 0 8952 0 1 -10
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_4  delaybuf0 $PDKPATH/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751558652
transform 1 0 888 0 1 -10
box -86 -86 1094 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_4  delaybuf1
timestamp 1751558652
transform 1 0 1896 0 1 -10
box -86 -86 1094 870
use gf180mcu_as_sc_mcu7t3v3__invz_2  delayen0
timestamp 1764933398
transform 1 0 7160 0 1 -10
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__invz_2  delayen1
timestamp 1764933398
transform 1 0 2904 0 1 -10
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__invz_2  delayenb1
timestamp 1764933398
transform 1 0 4920 0 1 -10
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  delayint0 $PDKPATH/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532043
transform 1 0 6712 0 1 -10
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fillcap_4  gf180mcu_as_sc_mcu7t3v3__fillcap_4_0 $PDKPATH/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532246
transform 1 0 10744 0 1 -10
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fillcap_4  gf180mcu_as_sc_mcu7t3v3__fillcap_4_1
timestamp 1751532246
transform 1 0 11192 0 1 -10
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fillcap_4  gf180mcu_as_sc_mcu7t3v3__fillcap_4_2
timestamp 1751532246
transform 1 0 -456 0 1 -10
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fillcap_4  gf180mcu_as_sc_mcu7t3v3__fillcap_4_3
timestamp 1751532246
transform 1 0 -904 0 1 -10
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  gf180mcu_as_sc_mcu7t3v3__diode_2_0 $PDKPATH/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532392
transform -1 0 -904 0 1 -10
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  gf180mcu_as_sc_mcu7t3v3__diode_2_1
timestamp 1751532392
transform -1 0 11864 0 1 -10
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  gf180mcu_as_sc_mcu7t3v3__tap_2_0 $PDKPATH/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1759751540
transform -1 0 12088 0 1 -10
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  gf180mcu_as_sc_mcu7t3v3__tap_2_1
timestamp 1759751540
transform -1 0 -1128 0 1 -10
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  gf180mcu_as_sc_mcu7t3v3__tap_2_2
timestamp 1759751540
transform 1 0 4696 0 1 -10
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  trim0bar
timestamp 1751532043
transform 1 0 -8 0 1 -10
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  trim1bar
timestamp 1751532043
transform 1 0 440 0 1 -10
box -86 -86 534 870
<< labels >>
flabel metal1 1760 304 1815 361 0 FreeSans 448 0 0 0 ts
flabel metal3 1090 466 1145 522 0 FreeSans 448 0 0 0 in
port 3 nsew
flabel metal1 -1128 714 -605 834 0 FreeSans 480 0 0 0 vdd
port 1 nsew
flabel metal1 -1128 -70 -605 50 0 FreeSans 480 0 0 0 vss
port 2 nsew
flabel metal3 -1326 18 -1271 74 0 FreeSans 448 0 0 0 trim[0]
port 4 nsew
flabel metal3 -1326 130 -1271 186 0 FreeSans 448 0 0 0 trim[1]
port 5 nsew
flabel metal3 6991 466 7045 522 0 FreeSans 480 0 0 0 d2
flabel metal3 8919 354 8977 410 0 FreeSans 448 0 0 0 out
port 6 nsew
flabel metal2 4216 632 4272 685 0 FreeSans 448 90 0 0 d1
flabel metal2 2592 633 2648 686 0 FreeSans 448 90 0 0 d0
<< end >>
