magic
tech gf180mcuD
magscale 1 10
timestamp 1765308861
<< nwell >>
rect 7000 607 7056 1270
<< metal1 >>
rect 374 2334 25324 2408
rect 374 2178 24655 2334
rect 24811 2178 25324 2334
rect 374 2108 25324 2178
rect 374 1478 17790 2108
rect 409 680 556 1478
rect 1397 1313 1443 1478
rect 1825 1309 1871 1478
rect 2258 1311 2304 1478
rect 2686 1311 2732 1478
rect 3064 923 3218 1478
rect 4908 1310 4954 1478
rect 5336 1311 5382 1478
rect 5764 1310 5810 1478
rect 6192 1310 6238 1478
rect 6358 933 6509 1478
rect 7361 704 7508 1478
rect 15845 874 17277 948
rect 15845 822 15967 874
rect 16019 822 16091 874
rect 16143 822 16215 874
rect 16267 822 16339 874
rect 16391 822 16463 874
rect 16515 822 16587 874
rect 16639 822 16711 874
rect 16763 822 16835 874
rect 16887 822 16959 874
rect 17011 822 17083 874
rect 17135 822 17277 874
rect 15845 750 17277 822
rect 15845 698 15967 750
rect 16019 698 16091 750
rect 16143 698 16215 750
rect 16267 698 16339 750
rect 16391 698 16463 750
rect 16515 698 16587 750
rect 16639 698 16711 750
rect 16763 698 16835 750
rect 16887 698 16959 750
rect 17011 698 17083 750
rect 17135 698 17277 750
rect 15845 626 17277 698
rect 15845 574 15967 626
rect 16019 574 16091 626
rect 16143 574 16215 626
rect 16267 574 16339 626
rect 16391 574 16463 626
rect 16515 574 16587 626
rect 16639 574 16711 626
rect 16763 574 16835 626
rect 16887 574 16959 626
rect 17011 574 17083 626
rect 17135 574 17277 626
rect 15845 502 17277 574
rect 7186 451 7580 473
rect 393 -357 505 381
rect 871 -357 1008 221
rect 1018 -357 1248 381
rect 3238 217 3468 381
rect 1607 -357 1653 -173
rect 2095 -357 2141 -176
rect 2583 -357 2629 -171
rect 3071 -357 3117 -171
rect 3238 -357 3601 217
rect 3977 -357 6761 381
rect 7186 295 7204 451
rect 7360 295 7580 451
rect 7186 273 7580 295
rect 15845 450 15967 502
rect 16019 450 16091 502
rect 16143 450 16215 502
rect 16267 450 16339 502
rect 16391 450 16463 502
rect 16515 450 16587 502
rect 16639 450 16711 502
rect 16763 450 16835 502
rect 16887 450 16959 502
rect 17011 450 17083 502
rect 17135 450 17277 502
rect 15845 378 17277 450
rect 15845 326 15967 378
rect 16019 326 16091 378
rect 16143 326 16215 378
rect 16267 326 16339 378
rect 16391 326 16463 378
rect 16515 326 16587 378
rect 16639 326 16711 378
rect 16763 326 16835 378
rect 16887 326 16959 378
rect 17011 326 17083 378
rect 17135 326 17277 378
rect 15845 254 17277 326
rect 15845 202 15967 254
rect 16019 202 16091 254
rect 16143 202 16215 254
rect 16267 202 16339 254
rect 16391 202 16463 254
rect 16515 202 16587 254
rect 16639 202 16711 254
rect 16763 202 16835 254
rect 16887 202 16959 254
rect 17011 202 17083 254
rect 17135 202 17277 254
rect 15845 130 17277 202
rect 15845 78 15967 130
rect 16019 78 16091 130
rect 16143 78 16215 130
rect 16267 78 16339 130
rect 16391 78 16463 130
rect 16515 78 16587 130
rect 16639 78 16711 130
rect 16763 78 16835 130
rect 16887 78 16959 130
rect 17011 78 17083 130
rect 17135 78 17277 130
rect 15845 6 17277 78
rect 15845 -46 15967 6
rect 16019 -46 16091 6
rect 16143 -46 16215 6
rect 16267 -46 16339 6
rect 16391 -46 16463 6
rect 16515 -46 16587 6
rect 16639 -46 16711 6
rect 16763 -46 16835 6
rect 16887 -46 16959 6
rect 17011 -46 17083 6
rect 17135 -46 17277 6
rect 15845 -118 17277 -46
rect 15845 -170 15967 -118
rect 16019 -170 16091 -118
rect 16143 -170 16215 -118
rect 16267 -170 16339 -118
rect 16391 -170 16463 -118
rect 16515 -170 16587 -118
rect 16639 -170 16711 -118
rect 16763 -170 16835 -118
rect 16887 -170 16959 -118
rect 17011 -170 17083 -118
rect 17135 -170 17277 -118
rect 15845 -242 17277 -170
rect 15845 -294 15967 -242
rect 16019 -294 16091 -242
rect 16143 -294 16215 -242
rect 16267 -294 16339 -242
rect 16391 -294 16463 -242
rect 16515 -294 16587 -242
rect 16639 -294 16711 -242
rect 16763 -294 16835 -242
rect 16887 -294 16959 -242
rect 17011 -294 17083 -242
rect 17135 -294 17277 -242
rect 15845 -357 17277 -294
rect 351 -366 25373 -357
rect 351 -418 15967 -366
rect 16019 -418 16091 -366
rect 16143 -418 16215 -366
rect 16267 -418 16339 -366
rect 16391 -418 16463 -366
rect 16515 -418 16587 -366
rect 16639 -418 16711 -366
rect 16763 -418 16835 -366
rect 16887 -418 16959 -366
rect 17011 -418 17083 -366
rect 17135 -418 25373 -366
rect 351 -657 25373 -418
rect 562 -825 758 -657
rect 837 -836 1320 -773
rect 1397 -836 1880 -773
rect 1957 -836 2440 -773
rect 2517 -779 3000 -773
rect 2517 -831 2684 -779
rect 2840 -831 3000 -779
rect 2517 -836 3000 -831
rect 3077 -836 3560 -773
rect 3637 -836 4120 -773
rect 4197 -836 4680 -773
rect 4757 -836 5240 -773
rect 5317 -836 5800 -773
rect 5877 -836 6360 -773
rect 6437 -836 6920 -773
rect 6997 -836 7480 -773
rect 7557 -836 8040 -773
rect 8117 -836 8600 -773
rect 8677 -836 9160 -773
rect 9237 -836 9720 -773
rect 9797 -836 10280 -773
rect 10357 -836 10840 -773
rect 10917 -836 11400 -773
rect 11477 -836 11960 -773
rect 12037 -836 12520 -773
rect 12597 -836 13080 -773
rect 13157 -836 13640 -773
rect 13717 -836 14200 -773
rect 14277 -836 14760 -773
rect 14837 -836 15320 -773
rect 15397 -836 15880 -773
rect 15957 -836 16440 -773
rect 16517 -836 17000 -773
rect 17077 -836 17560 -773
rect 17637 -836 18120 -773
rect 18197 -836 18680 -773
rect 18757 -836 19240 -773
rect 19317 -836 19800 -773
rect 19877 -836 20360 -773
rect 20437 -836 20920 -773
rect 20997 -836 21480 -773
rect 21557 -836 22040 -773
rect 22117 -836 22600 -773
rect 22677 -836 23160 -773
rect 23237 -836 23720 -773
rect 23797 -836 24280 -773
rect 24357 -836 24840 -773
rect 24917 -778 25124 -772
rect 24917 -830 24939 -778
rect 25095 -830 25124 -778
rect 24917 -833 25124 -830
rect 555 -6001 1038 -5938
rect 1115 -6001 1598 -5938
rect 1675 -6001 2158 -5938
rect 2235 -6001 2718 -5938
rect 2795 -6001 3278 -5938
rect 3355 -6001 3838 -5938
rect 3915 -6001 4398 -5938
rect 4475 -6001 4958 -5938
rect 5035 -6001 5518 -5938
rect 5595 -6001 6078 -5938
rect 6155 -6001 6638 -5938
rect 6715 -6001 7198 -5938
rect 7275 -6001 7758 -5938
rect 7835 -6001 8318 -5938
rect 8395 -6001 8878 -5938
rect 8955 -6001 9438 -5938
rect 9515 -6001 9998 -5938
rect 10075 -6001 10558 -5938
rect 10635 -6001 11118 -5938
rect 11195 -6001 11678 -5938
rect 11755 -6001 12238 -5938
rect 12315 -6001 12798 -5938
rect 12875 -6001 13358 -5938
rect 13435 -6001 13918 -5938
rect 13995 -6001 14478 -5938
rect 14555 -6001 15038 -5938
rect 15115 -6001 15598 -5938
rect 15675 -6001 16158 -5938
rect 16235 -6001 16718 -5938
rect 16795 -6001 17278 -5938
rect 17355 -6001 17838 -5938
rect 17915 -6001 18398 -5938
rect 18475 -6001 18958 -5938
rect 19035 -6001 19518 -5938
rect 19595 -6001 20078 -5938
rect 20155 -6001 20638 -5938
rect 20715 -6001 21198 -5938
rect 21275 -6001 21758 -5938
rect 21835 -6001 22318 -5938
rect 22395 -6001 22878 -5938
rect 22955 -6001 23438 -5938
rect 23515 -6001 23998 -5938
rect 24075 -6001 24558 -5938
rect 24635 -6001 25118 -5938
<< via1 >>
rect 24655 2178 24811 2334
rect 15967 822 16019 874
rect 16091 822 16143 874
rect 16215 822 16267 874
rect 16339 822 16391 874
rect 16463 822 16515 874
rect 16587 822 16639 874
rect 16711 822 16763 874
rect 16835 822 16887 874
rect 16959 822 17011 874
rect 17083 822 17135 874
rect 15967 698 16019 750
rect 16091 698 16143 750
rect 16215 698 16267 750
rect 16339 698 16391 750
rect 16463 698 16515 750
rect 16587 698 16639 750
rect 16711 698 16763 750
rect 16835 698 16887 750
rect 16959 698 17011 750
rect 17083 698 17135 750
rect 15967 574 16019 626
rect 16091 574 16143 626
rect 16215 574 16267 626
rect 16339 574 16391 626
rect 16463 574 16515 626
rect 16587 574 16639 626
rect 16711 574 16763 626
rect 16835 574 16887 626
rect 16959 574 17011 626
rect 17083 574 17135 626
rect 7204 295 7360 451
rect 15967 450 16019 502
rect 16091 450 16143 502
rect 16215 450 16267 502
rect 16339 450 16391 502
rect 16463 450 16515 502
rect 16587 450 16639 502
rect 16711 450 16763 502
rect 16835 450 16887 502
rect 16959 450 17011 502
rect 17083 450 17135 502
rect 15967 326 16019 378
rect 16091 326 16143 378
rect 16215 326 16267 378
rect 16339 326 16391 378
rect 16463 326 16515 378
rect 16587 326 16639 378
rect 16711 326 16763 378
rect 16835 326 16887 378
rect 16959 326 17011 378
rect 17083 326 17135 378
rect 15967 202 16019 254
rect 16091 202 16143 254
rect 16215 202 16267 254
rect 16339 202 16391 254
rect 16463 202 16515 254
rect 16587 202 16639 254
rect 16711 202 16763 254
rect 16835 202 16887 254
rect 16959 202 17011 254
rect 17083 202 17135 254
rect 15967 78 16019 130
rect 16091 78 16143 130
rect 16215 78 16267 130
rect 16339 78 16391 130
rect 16463 78 16515 130
rect 16587 78 16639 130
rect 16711 78 16763 130
rect 16835 78 16887 130
rect 16959 78 17011 130
rect 17083 78 17135 130
rect 15967 -46 16019 6
rect 16091 -46 16143 6
rect 16215 -46 16267 6
rect 16339 -46 16391 6
rect 16463 -46 16515 6
rect 16587 -46 16639 6
rect 16711 -46 16763 6
rect 16835 -46 16887 6
rect 16959 -46 17011 6
rect 17083 -46 17135 6
rect 15967 -170 16019 -118
rect 16091 -170 16143 -118
rect 16215 -170 16267 -118
rect 16339 -170 16391 -118
rect 16463 -170 16515 -118
rect 16587 -170 16639 -118
rect 16711 -170 16763 -118
rect 16835 -170 16887 -118
rect 16959 -170 17011 -118
rect 17083 -170 17135 -118
rect 15967 -294 16019 -242
rect 16091 -294 16143 -242
rect 16215 -294 16267 -242
rect 16339 -294 16391 -242
rect 16463 -294 16515 -242
rect 16587 -294 16639 -242
rect 16711 -294 16763 -242
rect 16835 -294 16887 -242
rect 16959 -294 17011 -242
rect 17083 -294 17135 -242
rect 15967 -418 16019 -366
rect 16091 -418 16143 -366
rect 16215 -418 16267 -366
rect 16339 -418 16391 -366
rect 16463 -418 16515 -366
rect 16587 -418 16639 -366
rect 16711 -418 16763 -366
rect 16835 -418 16887 -366
rect 16959 -418 17011 -366
rect 17083 -418 17135 -366
rect 2684 -831 2840 -779
rect 24939 -830 25095 -778
<< metal2 >>
rect 24594 2334 24869 2392
rect 24594 2178 24655 2334
rect 24811 2178 24869 2334
rect 24594 2127 24869 2178
rect 654 749 711 1267
rect 921 1004 2919 1206
rect 3432 1017 3716 1217
rect 1037 869 1093 1004
rect 804 749 860 849
rect 1037 813 3380 869
rect 3785 749 3841 825
rect 654 693 3841 749
rect 654 562 711 693
rect 3926 622 3982 1275
rect 607 505 711 562
rect 3296 566 3982 622
rect 4145 862 4203 1264
rect 4433 1027 5997 1208
rect 4145 806 4270 862
rect 4541 861 4602 1027
rect 6726 1023 7022 1218
rect 4145 739 4203 806
rect 4541 803 6672 861
rect 7091 739 7149 853
rect 4145 681 7149 739
rect 607 119 664 505
rect 3296 290 3352 566
rect 4145 507 4203 681
rect 3858 449 4203 507
rect 7220 473 7278 1272
rect 15845 876 17277 948
rect 15845 820 15965 876
rect 16021 820 16089 876
rect 16145 820 16213 876
rect 16269 820 16337 876
rect 16393 820 16461 876
rect 16517 820 16585 876
rect 16641 820 16709 876
rect 16765 820 16833 876
rect 16889 820 16957 876
rect 17013 820 17081 876
rect 17137 820 17277 876
rect 15845 752 17277 820
rect 15845 696 15965 752
rect 16021 696 16089 752
rect 16145 696 16213 752
rect 16269 696 16337 752
rect 16393 696 16461 752
rect 16517 696 16585 752
rect 16641 696 16709 752
rect 16765 696 16833 752
rect 16889 696 16957 752
rect 17013 696 17081 752
rect 17137 696 17277 752
rect 15845 628 17277 696
rect 15845 572 15965 628
rect 16021 572 16089 628
rect 16145 572 16213 628
rect 16269 572 16337 628
rect 16393 572 16461 628
rect 16517 572 16585 628
rect 16641 572 16709 628
rect 16765 572 16833 628
rect 16889 572 16957 628
rect 17013 572 17081 628
rect 17137 572 17277 628
rect 15845 504 17277 572
rect 7186 451 7633 473
rect 1437 222 3796 290
rect 3296 107 3352 222
rect 1393 -83 3352 107
rect 1393 -86 3341 -83
rect 3858 -195 3916 449
rect 7186 295 7204 451
rect 7360 295 7633 451
rect 7186 273 7633 295
rect 15845 448 15965 504
rect 16021 448 16089 504
rect 16145 448 16213 504
rect 16269 448 16337 504
rect 16393 448 16461 504
rect 16517 448 16585 504
rect 16641 448 16709 504
rect 16765 448 16833 504
rect 16889 448 16957 504
rect 17013 448 17081 504
rect 17137 448 17277 504
rect 15845 380 17277 448
rect 15845 324 15965 380
rect 16021 324 16089 380
rect 16145 324 16213 380
rect 16269 324 16337 380
rect 16393 324 16461 380
rect 16517 324 16585 380
rect 16641 324 16709 380
rect 16765 324 16833 380
rect 16889 324 16957 380
rect 17013 324 17081 380
rect 17137 324 17277 380
rect 15845 256 17277 324
rect 15845 200 15965 256
rect 16021 200 16089 256
rect 16145 200 16213 256
rect 16269 200 16337 256
rect 16393 200 16461 256
rect 16517 200 16585 256
rect 16641 200 16709 256
rect 16765 200 16833 256
rect 16889 200 16957 256
rect 17013 200 17081 256
rect 17137 200 17277 256
rect 15845 132 17277 200
rect 15845 76 15965 132
rect 16021 76 16089 132
rect 16145 76 16213 132
rect 16269 76 16337 132
rect 16393 76 16461 132
rect 16517 76 16585 132
rect 16641 76 16709 132
rect 16765 76 16833 132
rect 16889 76 16957 132
rect 17013 76 17081 132
rect 17137 76 17277 132
rect 15845 8 17277 76
rect 15845 -48 15965 8
rect 16021 -48 16089 8
rect 16145 -48 16213 8
rect 16269 -48 16337 8
rect 16393 -48 16461 8
rect 16517 -48 16585 8
rect 16641 -48 16709 8
rect 16765 -48 16833 8
rect 16889 -48 16957 8
rect 17013 -48 17081 8
rect 17137 -48 17277 8
rect 15845 -116 17277 -48
rect 15845 -172 15965 -116
rect 16021 -172 16089 -116
rect 16145 -172 16213 -116
rect 16269 -172 16337 -116
rect 16393 -172 16461 -116
rect 16517 -172 16585 -116
rect 16641 -172 16709 -116
rect 16765 -172 16833 -116
rect 16889 -172 16957 -116
rect 17013 -172 17081 -116
rect 17137 -172 17277 -116
rect 724 -510 787 -234
rect 15845 -240 17277 -172
rect 15845 -296 15965 -240
rect 16021 -296 16089 -240
rect 16145 -296 16213 -240
rect 16269 -296 16337 -240
rect 16393 -296 16461 -240
rect 16517 -296 16585 -240
rect 16641 -296 16709 -240
rect 16765 -296 16833 -240
rect 16889 -296 16957 -240
rect 17013 -296 17081 -240
rect 17137 -296 17277 -240
rect 15845 -364 17277 -296
rect 24641 -202 24800 2127
rect 24641 -361 25100 -202
rect 15845 -420 15965 -364
rect 16021 -420 16089 -364
rect 16145 -420 16213 -364
rect 16269 -420 16337 -364
rect 16393 -420 16461 -364
rect 16517 -420 16585 -364
rect 16641 -420 16709 -364
rect 16765 -420 16833 -364
rect 16889 -420 16957 -364
rect 17013 -420 17081 -364
rect 17137 -420 17277 -364
rect 15845 -500 17277 -420
rect 724 -573 2781 -510
rect 2718 -773 2781 -573
rect 24941 -772 25100 -361
rect 2624 -779 2903 -773
rect 2624 -831 2684 -779
rect 2840 -831 2903 -779
rect 2624 -835 2903 -831
rect 24916 -778 25123 -772
rect 24916 -830 24939 -778
rect 25095 -830 25123 -778
rect 24916 -834 25123 -830
<< via2 >>
rect 15965 874 16021 876
rect 15965 822 15967 874
rect 15967 822 16019 874
rect 16019 822 16021 874
rect 15965 820 16021 822
rect 16089 874 16145 876
rect 16089 822 16091 874
rect 16091 822 16143 874
rect 16143 822 16145 874
rect 16089 820 16145 822
rect 16213 874 16269 876
rect 16213 822 16215 874
rect 16215 822 16267 874
rect 16267 822 16269 874
rect 16213 820 16269 822
rect 16337 874 16393 876
rect 16337 822 16339 874
rect 16339 822 16391 874
rect 16391 822 16393 874
rect 16337 820 16393 822
rect 16461 874 16517 876
rect 16461 822 16463 874
rect 16463 822 16515 874
rect 16515 822 16517 874
rect 16461 820 16517 822
rect 16585 874 16641 876
rect 16585 822 16587 874
rect 16587 822 16639 874
rect 16639 822 16641 874
rect 16585 820 16641 822
rect 16709 874 16765 876
rect 16709 822 16711 874
rect 16711 822 16763 874
rect 16763 822 16765 874
rect 16709 820 16765 822
rect 16833 874 16889 876
rect 16833 822 16835 874
rect 16835 822 16887 874
rect 16887 822 16889 874
rect 16833 820 16889 822
rect 16957 874 17013 876
rect 16957 822 16959 874
rect 16959 822 17011 874
rect 17011 822 17013 874
rect 16957 820 17013 822
rect 17081 874 17137 876
rect 17081 822 17083 874
rect 17083 822 17135 874
rect 17135 822 17137 874
rect 17081 820 17137 822
rect 15965 750 16021 752
rect 15965 698 15967 750
rect 15967 698 16019 750
rect 16019 698 16021 750
rect 15965 696 16021 698
rect 16089 750 16145 752
rect 16089 698 16091 750
rect 16091 698 16143 750
rect 16143 698 16145 750
rect 16089 696 16145 698
rect 16213 750 16269 752
rect 16213 698 16215 750
rect 16215 698 16267 750
rect 16267 698 16269 750
rect 16213 696 16269 698
rect 16337 750 16393 752
rect 16337 698 16339 750
rect 16339 698 16391 750
rect 16391 698 16393 750
rect 16337 696 16393 698
rect 16461 750 16517 752
rect 16461 698 16463 750
rect 16463 698 16515 750
rect 16515 698 16517 750
rect 16461 696 16517 698
rect 16585 750 16641 752
rect 16585 698 16587 750
rect 16587 698 16639 750
rect 16639 698 16641 750
rect 16585 696 16641 698
rect 16709 750 16765 752
rect 16709 698 16711 750
rect 16711 698 16763 750
rect 16763 698 16765 750
rect 16709 696 16765 698
rect 16833 750 16889 752
rect 16833 698 16835 750
rect 16835 698 16887 750
rect 16887 698 16889 750
rect 16833 696 16889 698
rect 16957 750 17013 752
rect 16957 698 16959 750
rect 16959 698 17011 750
rect 17011 698 17013 750
rect 16957 696 17013 698
rect 17081 750 17137 752
rect 17081 698 17083 750
rect 17083 698 17135 750
rect 17135 698 17137 750
rect 17081 696 17137 698
rect 15965 626 16021 628
rect 15965 574 15967 626
rect 15967 574 16019 626
rect 16019 574 16021 626
rect 15965 572 16021 574
rect 16089 626 16145 628
rect 16089 574 16091 626
rect 16091 574 16143 626
rect 16143 574 16145 626
rect 16089 572 16145 574
rect 16213 626 16269 628
rect 16213 574 16215 626
rect 16215 574 16267 626
rect 16267 574 16269 626
rect 16213 572 16269 574
rect 16337 626 16393 628
rect 16337 574 16339 626
rect 16339 574 16391 626
rect 16391 574 16393 626
rect 16337 572 16393 574
rect 16461 626 16517 628
rect 16461 574 16463 626
rect 16463 574 16515 626
rect 16515 574 16517 626
rect 16461 572 16517 574
rect 16585 626 16641 628
rect 16585 574 16587 626
rect 16587 574 16639 626
rect 16639 574 16641 626
rect 16585 572 16641 574
rect 16709 626 16765 628
rect 16709 574 16711 626
rect 16711 574 16763 626
rect 16763 574 16765 626
rect 16709 572 16765 574
rect 16833 626 16889 628
rect 16833 574 16835 626
rect 16835 574 16887 626
rect 16887 574 16889 626
rect 16833 572 16889 574
rect 16957 626 17013 628
rect 16957 574 16959 626
rect 16959 574 17011 626
rect 17011 574 17013 626
rect 16957 572 17013 574
rect 17081 626 17137 628
rect 17081 574 17083 626
rect 17083 574 17135 626
rect 17135 574 17137 626
rect 17081 572 17137 574
rect 15965 502 16021 504
rect 15965 450 15967 502
rect 15967 450 16019 502
rect 16019 450 16021 502
rect 15965 448 16021 450
rect 16089 502 16145 504
rect 16089 450 16091 502
rect 16091 450 16143 502
rect 16143 450 16145 502
rect 16089 448 16145 450
rect 16213 502 16269 504
rect 16213 450 16215 502
rect 16215 450 16267 502
rect 16267 450 16269 502
rect 16213 448 16269 450
rect 16337 502 16393 504
rect 16337 450 16339 502
rect 16339 450 16391 502
rect 16391 450 16393 502
rect 16337 448 16393 450
rect 16461 502 16517 504
rect 16461 450 16463 502
rect 16463 450 16515 502
rect 16515 450 16517 502
rect 16461 448 16517 450
rect 16585 502 16641 504
rect 16585 450 16587 502
rect 16587 450 16639 502
rect 16639 450 16641 502
rect 16585 448 16641 450
rect 16709 502 16765 504
rect 16709 450 16711 502
rect 16711 450 16763 502
rect 16763 450 16765 502
rect 16709 448 16765 450
rect 16833 502 16889 504
rect 16833 450 16835 502
rect 16835 450 16887 502
rect 16887 450 16889 502
rect 16833 448 16889 450
rect 16957 502 17013 504
rect 16957 450 16959 502
rect 16959 450 17011 502
rect 17011 450 17013 502
rect 16957 448 17013 450
rect 17081 502 17137 504
rect 17081 450 17083 502
rect 17083 450 17135 502
rect 17135 450 17137 502
rect 17081 448 17137 450
rect 15965 378 16021 380
rect 15965 326 15967 378
rect 15967 326 16019 378
rect 16019 326 16021 378
rect 15965 324 16021 326
rect 16089 378 16145 380
rect 16089 326 16091 378
rect 16091 326 16143 378
rect 16143 326 16145 378
rect 16089 324 16145 326
rect 16213 378 16269 380
rect 16213 326 16215 378
rect 16215 326 16267 378
rect 16267 326 16269 378
rect 16213 324 16269 326
rect 16337 378 16393 380
rect 16337 326 16339 378
rect 16339 326 16391 378
rect 16391 326 16393 378
rect 16337 324 16393 326
rect 16461 378 16517 380
rect 16461 326 16463 378
rect 16463 326 16515 378
rect 16515 326 16517 378
rect 16461 324 16517 326
rect 16585 378 16641 380
rect 16585 326 16587 378
rect 16587 326 16639 378
rect 16639 326 16641 378
rect 16585 324 16641 326
rect 16709 378 16765 380
rect 16709 326 16711 378
rect 16711 326 16763 378
rect 16763 326 16765 378
rect 16709 324 16765 326
rect 16833 378 16889 380
rect 16833 326 16835 378
rect 16835 326 16887 378
rect 16887 326 16889 378
rect 16833 324 16889 326
rect 16957 378 17013 380
rect 16957 326 16959 378
rect 16959 326 17011 378
rect 17011 326 17013 378
rect 16957 324 17013 326
rect 17081 378 17137 380
rect 17081 326 17083 378
rect 17083 326 17135 378
rect 17135 326 17137 378
rect 17081 324 17137 326
rect 15965 254 16021 256
rect 15965 202 15967 254
rect 15967 202 16019 254
rect 16019 202 16021 254
rect 15965 200 16021 202
rect 16089 254 16145 256
rect 16089 202 16091 254
rect 16091 202 16143 254
rect 16143 202 16145 254
rect 16089 200 16145 202
rect 16213 254 16269 256
rect 16213 202 16215 254
rect 16215 202 16267 254
rect 16267 202 16269 254
rect 16213 200 16269 202
rect 16337 254 16393 256
rect 16337 202 16339 254
rect 16339 202 16391 254
rect 16391 202 16393 254
rect 16337 200 16393 202
rect 16461 254 16517 256
rect 16461 202 16463 254
rect 16463 202 16515 254
rect 16515 202 16517 254
rect 16461 200 16517 202
rect 16585 254 16641 256
rect 16585 202 16587 254
rect 16587 202 16639 254
rect 16639 202 16641 254
rect 16585 200 16641 202
rect 16709 254 16765 256
rect 16709 202 16711 254
rect 16711 202 16763 254
rect 16763 202 16765 254
rect 16709 200 16765 202
rect 16833 254 16889 256
rect 16833 202 16835 254
rect 16835 202 16887 254
rect 16887 202 16889 254
rect 16833 200 16889 202
rect 16957 254 17013 256
rect 16957 202 16959 254
rect 16959 202 17011 254
rect 17011 202 17013 254
rect 16957 200 17013 202
rect 17081 254 17137 256
rect 17081 202 17083 254
rect 17083 202 17135 254
rect 17135 202 17137 254
rect 17081 200 17137 202
rect 15965 130 16021 132
rect 15965 78 15967 130
rect 15967 78 16019 130
rect 16019 78 16021 130
rect 15965 76 16021 78
rect 16089 130 16145 132
rect 16089 78 16091 130
rect 16091 78 16143 130
rect 16143 78 16145 130
rect 16089 76 16145 78
rect 16213 130 16269 132
rect 16213 78 16215 130
rect 16215 78 16267 130
rect 16267 78 16269 130
rect 16213 76 16269 78
rect 16337 130 16393 132
rect 16337 78 16339 130
rect 16339 78 16391 130
rect 16391 78 16393 130
rect 16337 76 16393 78
rect 16461 130 16517 132
rect 16461 78 16463 130
rect 16463 78 16515 130
rect 16515 78 16517 130
rect 16461 76 16517 78
rect 16585 130 16641 132
rect 16585 78 16587 130
rect 16587 78 16639 130
rect 16639 78 16641 130
rect 16585 76 16641 78
rect 16709 130 16765 132
rect 16709 78 16711 130
rect 16711 78 16763 130
rect 16763 78 16765 130
rect 16709 76 16765 78
rect 16833 130 16889 132
rect 16833 78 16835 130
rect 16835 78 16887 130
rect 16887 78 16889 130
rect 16833 76 16889 78
rect 16957 130 17013 132
rect 16957 78 16959 130
rect 16959 78 17011 130
rect 17011 78 17013 130
rect 16957 76 17013 78
rect 17081 130 17137 132
rect 17081 78 17083 130
rect 17083 78 17135 130
rect 17135 78 17137 130
rect 17081 76 17137 78
rect 15965 6 16021 8
rect 15965 -46 15967 6
rect 15967 -46 16019 6
rect 16019 -46 16021 6
rect 15965 -48 16021 -46
rect 16089 6 16145 8
rect 16089 -46 16091 6
rect 16091 -46 16143 6
rect 16143 -46 16145 6
rect 16089 -48 16145 -46
rect 16213 6 16269 8
rect 16213 -46 16215 6
rect 16215 -46 16267 6
rect 16267 -46 16269 6
rect 16213 -48 16269 -46
rect 16337 6 16393 8
rect 16337 -46 16339 6
rect 16339 -46 16391 6
rect 16391 -46 16393 6
rect 16337 -48 16393 -46
rect 16461 6 16517 8
rect 16461 -46 16463 6
rect 16463 -46 16515 6
rect 16515 -46 16517 6
rect 16461 -48 16517 -46
rect 16585 6 16641 8
rect 16585 -46 16587 6
rect 16587 -46 16639 6
rect 16639 -46 16641 6
rect 16585 -48 16641 -46
rect 16709 6 16765 8
rect 16709 -46 16711 6
rect 16711 -46 16763 6
rect 16763 -46 16765 6
rect 16709 -48 16765 -46
rect 16833 6 16889 8
rect 16833 -46 16835 6
rect 16835 -46 16887 6
rect 16887 -46 16889 6
rect 16833 -48 16889 -46
rect 16957 6 17013 8
rect 16957 -46 16959 6
rect 16959 -46 17011 6
rect 17011 -46 17013 6
rect 16957 -48 17013 -46
rect 17081 6 17137 8
rect 17081 -46 17083 6
rect 17083 -46 17135 6
rect 17135 -46 17137 6
rect 17081 -48 17137 -46
rect 15965 -118 16021 -116
rect 15965 -170 15967 -118
rect 15967 -170 16019 -118
rect 16019 -170 16021 -118
rect 15965 -172 16021 -170
rect 16089 -118 16145 -116
rect 16089 -170 16091 -118
rect 16091 -170 16143 -118
rect 16143 -170 16145 -118
rect 16089 -172 16145 -170
rect 16213 -118 16269 -116
rect 16213 -170 16215 -118
rect 16215 -170 16267 -118
rect 16267 -170 16269 -118
rect 16213 -172 16269 -170
rect 16337 -118 16393 -116
rect 16337 -170 16339 -118
rect 16339 -170 16391 -118
rect 16391 -170 16393 -118
rect 16337 -172 16393 -170
rect 16461 -118 16517 -116
rect 16461 -170 16463 -118
rect 16463 -170 16515 -118
rect 16515 -170 16517 -118
rect 16461 -172 16517 -170
rect 16585 -118 16641 -116
rect 16585 -170 16587 -118
rect 16587 -170 16639 -118
rect 16639 -170 16641 -118
rect 16585 -172 16641 -170
rect 16709 -118 16765 -116
rect 16709 -170 16711 -118
rect 16711 -170 16763 -118
rect 16763 -170 16765 -118
rect 16709 -172 16765 -170
rect 16833 -118 16889 -116
rect 16833 -170 16835 -118
rect 16835 -170 16887 -118
rect 16887 -170 16889 -118
rect 16833 -172 16889 -170
rect 16957 -118 17013 -116
rect 16957 -170 16959 -118
rect 16959 -170 17011 -118
rect 17011 -170 17013 -118
rect 16957 -172 17013 -170
rect 17081 -118 17137 -116
rect 17081 -170 17083 -118
rect 17083 -170 17135 -118
rect 17135 -170 17137 -118
rect 17081 -172 17137 -170
rect 15965 -242 16021 -240
rect 15965 -294 15967 -242
rect 15967 -294 16019 -242
rect 16019 -294 16021 -242
rect 15965 -296 16021 -294
rect 16089 -242 16145 -240
rect 16089 -294 16091 -242
rect 16091 -294 16143 -242
rect 16143 -294 16145 -242
rect 16089 -296 16145 -294
rect 16213 -242 16269 -240
rect 16213 -294 16215 -242
rect 16215 -294 16267 -242
rect 16267 -294 16269 -242
rect 16213 -296 16269 -294
rect 16337 -242 16393 -240
rect 16337 -294 16339 -242
rect 16339 -294 16391 -242
rect 16391 -294 16393 -242
rect 16337 -296 16393 -294
rect 16461 -242 16517 -240
rect 16461 -294 16463 -242
rect 16463 -294 16515 -242
rect 16515 -294 16517 -242
rect 16461 -296 16517 -294
rect 16585 -242 16641 -240
rect 16585 -294 16587 -242
rect 16587 -294 16639 -242
rect 16639 -294 16641 -242
rect 16585 -296 16641 -294
rect 16709 -242 16765 -240
rect 16709 -294 16711 -242
rect 16711 -294 16763 -242
rect 16763 -294 16765 -242
rect 16709 -296 16765 -294
rect 16833 -242 16889 -240
rect 16833 -294 16835 -242
rect 16835 -294 16887 -242
rect 16887 -294 16889 -242
rect 16833 -296 16889 -294
rect 16957 -242 17013 -240
rect 16957 -294 16959 -242
rect 16959 -294 17011 -242
rect 17011 -294 17013 -242
rect 16957 -296 17013 -294
rect 17081 -242 17137 -240
rect 17081 -294 17083 -242
rect 17083 -294 17135 -242
rect 17135 -294 17137 -242
rect 17081 -296 17137 -294
rect 15965 -366 16021 -364
rect 15965 -418 15967 -366
rect 15967 -418 16019 -366
rect 16019 -418 16021 -366
rect 15965 -420 16021 -418
rect 16089 -366 16145 -364
rect 16089 -418 16091 -366
rect 16091 -418 16143 -366
rect 16143 -418 16145 -366
rect 16089 -420 16145 -418
rect 16213 -366 16269 -364
rect 16213 -418 16215 -366
rect 16215 -418 16267 -366
rect 16267 -418 16269 -366
rect 16213 -420 16269 -418
rect 16337 -366 16393 -364
rect 16337 -418 16339 -366
rect 16339 -418 16391 -366
rect 16391 -418 16393 -366
rect 16337 -420 16393 -418
rect 16461 -366 16517 -364
rect 16461 -418 16463 -366
rect 16463 -418 16515 -366
rect 16515 -418 16517 -366
rect 16461 -420 16517 -418
rect 16585 -366 16641 -364
rect 16585 -418 16587 -366
rect 16587 -418 16639 -366
rect 16639 -418 16641 -366
rect 16585 -420 16641 -418
rect 16709 -366 16765 -364
rect 16709 -418 16711 -366
rect 16711 -418 16763 -366
rect 16763 -418 16765 -366
rect 16709 -420 16765 -418
rect 16833 -366 16889 -364
rect 16833 -418 16835 -366
rect 16835 -418 16887 -366
rect 16887 -418 16889 -366
rect 16833 -420 16889 -418
rect 16957 -366 17013 -364
rect 16957 -418 16959 -366
rect 16959 -418 17011 -366
rect 17011 -418 17013 -366
rect 16957 -420 17013 -418
rect 17081 -366 17137 -364
rect 17081 -418 17083 -366
rect 17083 -418 17135 -366
rect 17135 -418 17137 -366
rect 17081 -420 17137 -418
<< metal3 >>
rect 15845 876 17277 948
rect 15845 820 15965 876
rect 16063 820 16089 876
rect 16187 820 16213 876
rect 16311 820 16337 876
rect 16435 820 16461 876
rect 16559 820 16585 876
rect 16683 820 16709 876
rect 16807 820 16833 876
rect 16931 820 16957 876
rect 17055 820 17081 876
rect 17179 820 17277 876
rect 15845 752 17277 820
rect 15845 696 15965 752
rect 16063 696 16089 752
rect 16187 696 16213 752
rect 16311 696 16337 752
rect 16435 696 16461 752
rect 16559 696 16585 752
rect 16683 696 16709 752
rect 16807 696 16833 752
rect 16931 696 16957 752
rect 17055 696 17081 752
rect 17179 696 17277 752
rect 15845 628 17277 696
rect 15845 572 15965 628
rect 16063 572 16089 628
rect 16187 572 16213 628
rect 16311 572 16337 628
rect 16435 572 16461 628
rect 16559 572 16585 628
rect 16683 572 16709 628
rect 16807 572 16833 628
rect 16931 572 16957 628
rect 17055 572 17081 628
rect 17179 572 17277 628
rect 15845 504 17277 572
rect 15845 448 15965 504
rect 16063 448 16089 504
rect 16187 448 16213 504
rect 16311 448 16337 504
rect 16435 448 16461 504
rect 16559 448 16585 504
rect 16683 448 16709 504
rect 16807 448 16833 504
rect 16931 448 16957 504
rect 17055 448 17081 504
rect 17179 448 17277 504
rect 15845 380 17277 448
rect 15845 324 15965 380
rect 16063 324 16089 380
rect 16187 324 16213 380
rect 16311 324 16337 380
rect 16435 324 16461 380
rect 16559 324 16585 380
rect 16683 324 16709 380
rect 16807 324 16833 380
rect 16931 324 16957 380
rect 17055 324 17081 380
rect 17179 324 17277 380
rect 15845 256 17277 324
rect 15845 200 15965 256
rect 16063 200 16089 256
rect 16187 200 16213 256
rect 16311 200 16337 256
rect 16435 200 16461 256
rect 16559 200 16585 256
rect 16683 200 16709 256
rect 16807 200 16833 256
rect 16931 200 16957 256
rect 17055 200 17081 256
rect 17179 200 17277 256
rect 15845 132 17277 200
rect 15845 76 15965 132
rect 16063 76 16089 132
rect 16187 76 16213 132
rect 16311 76 16337 132
rect 16435 76 16461 132
rect 16559 76 16585 132
rect 16683 76 16709 132
rect 16807 76 16833 132
rect 16931 76 16957 132
rect 17055 76 17081 132
rect 17179 76 17277 132
rect 15845 8 17277 76
rect 15845 -48 15965 8
rect 16063 -48 16089 8
rect 16187 -48 16213 8
rect 16311 -48 16337 8
rect 16435 -48 16461 8
rect 16559 -48 16585 8
rect 16683 -48 16709 8
rect 16807 -48 16833 8
rect 16931 -48 16957 8
rect 17055 -48 17081 8
rect 17179 -48 17277 8
rect 15845 -116 17277 -48
rect 15845 -172 15965 -116
rect 16063 -172 16089 -116
rect 16187 -172 16213 -116
rect 16311 -172 16337 -116
rect 16435 -172 16461 -116
rect 16559 -172 16585 -116
rect 16683 -172 16709 -116
rect 16807 -172 16833 -116
rect 16931 -172 16957 -116
rect 17055 -172 17081 -116
rect 17179 -172 17277 -116
rect 15845 -240 17277 -172
rect 15845 -296 15965 -240
rect 16063 -296 16089 -240
rect 16187 -296 16213 -240
rect 16311 -296 16337 -240
rect 16435 -296 16461 -240
rect 16559 -296 16585 -240
rect 16683 -296 16709 -240
rect 16807 -296 16833 -240
rect 16931 -296 16957 -240
rect 17055 -296 17081 -240
rect 17179 -296 17277 -240
rect 15845 -364 17277 -296
rect 15845 -420 15965 -364
rect 16063 -420 16089 -364
rect 16187 -420 16213 -364
rect 16311 -420 16337 -364
rect 16435 -420 16461 -364
rect 16559 -420 16585 -364
rect 16683 -420 16709 -364
rect 16807 -420 16833 -364
rect 16931 -420 16957 -364
rect 17055 -420 17081 -364
rect 17179 -420 17277 -364
rect 15845 -500 17277 -420
<< via3 >>
rect 16007 820 16021 876
rect 16021 820 16063 876
rect 16131 820 16145 876
rect 16145 820 16187 876
rect 16255 820 16269 876
rect 16269 820 16311 876
rect 16379 820 16393 876
rect 16393 820 16435 876
rect 16503 820 16517 876
rect 16517 820 16559 876
rect 16627 820 16641 876
rect 16641 820 16683 876
rect 16751 820 16765 876
rect 16765 820 16807 876
rect 16875 820 16889 876
rect 16889 820 16931 876
rect 16999 820 17013 876
rect 17013 820 17055 876
rect 17123 820 17137 876
rect 17137 820 17179 876
rect 16007 696 16021 752
rect 16021 696 16063 752
rect 16131 696 16145 752
rect 16145 696 16187 752
rect 16255 696 16269 752
rect 16269 696 16311 752
rect 16379 696 16393 752
rect 16393 696 16435 752
rect 16503 696 16517 752
rect 16517 696 16559 752
rect 16627 696 16641 752
rect 16641 696 16683 752
rect 16751 696 16765 752
rect 16765 696 16807 752
rect 16875 696 16889 752
rect 16889 696 16931 752
rect 16999 696 17013 752
rect 17013 696 17055 752
rect 17123 696 17137 752
rect 17137 696 17179 752
rect 16007 572 16021 628
rect 16021 572 16063 628
rect 16131 572 16145 628
rect 16145 572 16187 628
rect 16255 572 16269 628
rect 16269 572 16311 628
rect 16379 572 16393 628
rect 16393 572 16435 628
rect 16503 572 16517 628
rect 16517 572 16559 628
rect 16627 572 16641 628
rect 16641 572 16683 628
rect 16751 572 16765 628
rect 16765 572 16807 628
rect 16875 572 16889 628
rect 16889 572 16931 628
rect 16999 572 17013 628
rect 17013 572 17055 628
rect 17123 572 17137 628
rect 17137 572 17179 628
rect 16007 448 16021 504
rect 16021 448 16063 504
rect 16131 448 16145 504
rect 16145 448 16187 504
rect 16255 448 16269 504
rect 16269 448 16311 504
rect 16379 448 16393 504
rect 16393 448 16435 504
rect 16503 448 16517 504
rect 16517 448 16559 504
rect 16627 448 16641 504
rect 16641 448 16683 504
rect 16751 448 16765 504
rect 16765 448 16807 504
rect 16875 448 16889 504
rect 16889 448 16931 504
rect 16999 448 17013 504
rect 17013 448 17055 504
rect 17123 448 17137 504
rect 17137 448 17179 504
rect 16007 324 16021 380
rect 16021 324 16063 380
rect 16131 324 16145 380
rect 16145 324 16187 380
rect 16255 324 16269 380
rect 16269 324 16311 380
rect 16379 324 16393 380
rect 16393 324 16435 380
rect 16503 324 16517 380
rect 16517 324 16559 380
rect 16627 324 16641 380
rect 16641 324 16683 380
rect 16751 324 16765 380
rect 16765 324 16807 380
rect 16875 324 16889 380
rect 16889 324 16931 380
rect 16999 324 17013 380
rect 17013 324 17055 380
rect 17123 324 17137 380
rect 17137 324 17179 380
rect 16007 200 16021 256
rect 16021 200 16063 256
rect 16131 200 16145 256
rect 16145 200 16187 256
rect 16255 200 16269 256
rect 16269 200 16311 256
rect 16379 200 16393 256
rect 16393 200 16435 256
rect 16503 200 16517 256
rect 16517 200 16559 256
rect 16627 200 16641 256
rect 16641 200 16683 256
rect 16751 200 16765 256
rect 16765 200 16807 256
rect 16875 200 16889 256
rect 16889 200 16931 256
rect 16999 200 17013 256
rect 17013 200 17055 256
rect 17123 200 17137 256
rect 17137 200 17179 256
rect 16007 76 16021 132
rect 16021 76 16063 132
rect 16131 76 16145 132
rect 16145 76 16187 132
rect 16255 76 16269 132
rect 16269 76 16311 132
rect 16379 76 16393 132
rect 16393 76 16435 132
rect 16503 76 16517 132
rect 16517 76 16559 132
rect 16627 76 16641 132
rect 16641 76 16683 132
rect 16751 76 16765 132
rect 16765 76 16807 132
rect 16875 76 16889 132
rect 16889 76 16931 132
rect 16999 76 17013 132
rect 17013 76 17055 132
rect 17123 76 17137 132
rect 17137 76 17179 132
rect 16007 -48 16021 8
rect 16021 -48 16063 8
rect 16131 -48 16145 8
rect 16145 -48 16187 8
rect 16255 -48 16269 8
rect 16269 -48 16311 8
rect 16379 -48 16393 8
rect 16393 -48 16435 8
rect 16503 -48 16517 8
rect 16517 -48 16559 8
rect 16627 -48 16641 8
rect 16641 -48 16683 8
rect 16751 -48 16765 8
rect 16765 -48 16807 8
rect 16875 -48 16889 8
rect 16889 -48 16931 8
rect 16999 -48 17013 8
rect 17013 -48 17055 8
rect 17123 -48 17137 8
rect 17137 -48 17179 8
rect 16007 -172 16021 -116
rect 16021 -172 16063 -116
rect 16131 -172 16145 -116
rect 16145 -172 16187 -116
rect 16255 -172 16269 -116
rect 16269 -172 16311 -116
rect 16379 -172 16393 -116
rect 16393 -172 16435 -116
rect 16503 -172 16517 -116
rect 16517 -172 16559 -116
rect 16627 -172 16641 -116
rect 16641 -172 16683 -116
rect 16751 -172 16765 -116
rect 16765 -172 16807 -116
rect 16875 -172 16889 -116
rect 16889 -172 16931 -116
rect 16999 -172 17013 -116
rect 17013 -172 17055 -116
rect 17123 -172 17137 -116
rect 17137 -172 17179 -116
rect 16007 -296 16021 -240
rect 16021 -296 16063 -240
rect 16131 -296 16145 -240
rect 16145 -296 16187 -240
rect 16255 -296 16269 -240
rect 16269 -296 16311 -240
rect 16379 -296 16393 -240
rect 16393 -296 16435 -240
rect 16503 -296 16517 -240
rect 16517 -296 16559 -240
rect 16627 -296 16641 -240
rect 16641 -296 16683 -240
rect 16751 -296 16765 -240
rect 16765 -296 16807 -240
rect 16875 -296 16889 -240
rect 16889 -296 16931 -240
rect 16999 -296 17013 -240
rect 17013 -296 17055 -240
rect 17123 -296 17137 -240
rect 17137 -296 17179 -240
rect 16007 -420 16021 -364
rect 16021 -420 16063 -364
rect 16131 -420 16145 -364
rect 16145 -420 16187 -364
rect 16255 -420 16269 -364
rect 16269 -420 16311 -364
rect 16379 -420 16393 -364
rect 16393 -420 16435 -364
rect 16503 -420 16517 -364
rect 16517 -420 16559 -364
rect 16627 -420 16641 -364
rect 16641 -420 16683 -364
rect 16751 -420 16765 -364
rect 16765 -420 16807 -364
rect 16875 -420 16889 -364
rect 16889 -420 16931 -364
rect 16999 -420 17013 -364
rect 17013 -420 17055 -364
rect 17123 -420 17137 -364
rect 17137 -420 17179 -364
<< metal4 >>
rect 15955 876 17277 948
rect 15955 820 16007 876
rect 16063 820 16131 876
rect 16187 820 16255 876
rect 16311 820 16379 876
rect 16435 820 16503 876
rect 16559 820 16627 876
rect 16683 820 16751 876
rect 16807 820 16875 876
rect 16931 820 16999 876
rect 17055 820 17123 876
rect 17179 820 17277 876
rect 15955 752 17277 820
rect 15955 696 16007 752
rect 16063 696 16131 752
rect 16187 696 16255 752
rect 16311 696 16379 752
rect 16435 696 16503 752
rect 16559 696 16627 752
rect 16683 696 16751 752
rect 16807 696 16875 752
rect 16931 696 16999 752
rect 17055 696 17123 752
rect 17179 696 17277 752
rect 15955 628 17277 696
rect 15955 572 16007 628
rect 16063 572 16131 628
rect 16187 572 16255 628
rect 16311 572 16379 628
rect 16435 572 16503 628
rect 16559 572 16627 628
rect 16683 572 16751 628
rect 16807 572 16875 628
rect 16931 572 16999 628
rect 17055 572 17123 628
rect 17179 572 17277 628
rect 15955 504 17277 572
rect 15955 448 16007 504
rect 16063 448 16131 504
rect 16187 448 16255 504
rect 16311 448 16379 504
rect 16435 448 16503 504
rect 16559 448 16627 504
rect 16683 448 16751 504
rect 16807 448 16875 504
rect 16931 448 16999 504
rect 17055 448 17123 504
rect 17179 448 17277 504
rect 15955 380 17277 448
rect 15955 324 16007 380
rect 16063 324 16131 380
rect 16187 324 16255 380
rect 16311 324 16379 380
rect 16435 324 16503 380
rect 16559 324 16627 380
rect 16683 324 16751 380
rect 16807 324 16875 380
rect 16931 324 16999 380
rect 17055 324 17123 380
rect 17179 324 17277 380
rect 15955 256 17277 324
rect 15955 200 16007 256
rect 16063 200 16131 256
rect 16187 200 16255 256
rect 16311 200 16379 256
rect 16435 200 16503 256
rect 16559 200 16627 256
rect 16683 200 16751 256
rect 16807 200 16875 256
rect 16931 200 16999 256
rect 17055 200 17123 256
rect 17179 200 17277 256
rect 15955 132 17277 200
rect 15955 76 16007 132
rect 16063 76 16131 132
rect 16187 76 16255 132
rect 16311 76 16379 132
rect 16435 76 16503 132
rect 16559 76 16627 132
rect 16683 76 16751 132
rect 16807 76 16875 132
rect 16931 76 16999 132
rect 17055 76 17123 132
rect 17179 76 17277 132
rect 15955 8 17277 76
rect 15955 -48 16007 8
rect 16063 -48 16131 8
rect 16187 -48 16255 8
rect 16311 -48 16379 8
rect 16435 -48 16503 8
rect 16559 -48 16627 8
rect 16683 -48 16751 8
rect 16807 -48 16875 8
rect 16931 -48 16999 8
rect 17055 -48 17123 8
rect 17179 -48 17277 8
rect 15955 -116 17277 -48
rect 15955 -172 16007 -116
rect 16063 -172 16131 -116
rect 16187 -172 16255 -116
rect 16311 -172 16379 -116
rect 16435 -172 16503 -116
rect 16559 -172 16627 -116
rect 16683 -172 16751 -116
rect 16807 -172 16875 -116
rect 16931 -172 16999 -116
rect 17055 -172 17123 -116
rect 17179 -172 17277 -116
rect 15955 -240 17277 -172
rect 15955 -296 16007 -240
rect 16063 -296 16131 -240
rect 16187 -296 16255 -240
rect 16311 -296 16379 -240
rect 16435 -296 16503 -240
rect 16559 -296 16627 -240
rect 16683 -296 16751 -240
rect 16807 -296 16875 -240
rect 16931 -296 16999 -240
rect 17055 -296 17123 -240
rect 17179 -296 17277 -240
rect 15955 -364 17277 -296
rect 15955 -420 16007 -364
rect 16063 -420 16131 -364
rect 16187 -420 16255 -364
rect 16311 -420 16379 -364
rect 16435 -420 16503 -364
rect 16559 -420 16627 -364
rect 16683 -420 16751 -364
rect 16807 -420 16875 -364
rect 16931 -420 16999 -364
rect 17055 -420 17123 -364
rect 17179 -420 17277 -364
rect 15955 -500 17277 -420
use nmos_6p0_BJPB5U  nmos_6p0_BJPB5U_0
timestamp 1765308861
transform 1 0 3722 0 1 -4
box -334 -432 334 432
use nmos_6p0_BJXXPT  nmos_6p0_BJXXPT_0
timestamp 1765308861
transform 1 0 2242 0 1 8
box -1066 -432 1066 432
use pmos_6p0_CYEQN4  pmos_6p0_CYEQN4_0
timestamp 1765308861
transform 1 0 7107 0 1 1093
box -368 -486 378 486
use pmos_6p0_EYEQQM  pmos_6p0_EYEQQM_0
timestamp 1765308861
transform 1 0 5501 0 1 1093
box -1050 -486 980 486
use pmos_6p0_HUEQQM  pmos_6p0_HUEQQM_0
timestamp 1765308861
transform 1 0 2068 0 1 1093
box -1128 -486 1121 486
use ppolyf_u_1k_6p0_TRTT7C  ppolyf_u_1k_6p0_TRTT7C_0
timestamp 1765308861
transform 1 0 12839 0 1 -3388
box -12578 -2920 12578 2920
use via_cont_0p6um  via_cont_0p6um_0
timestamp 1765308861
transform 1 0 724 0 1 -55
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_1
timestamp 1765308861
transform 1 0 1483 0 1 432
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_2
timestamp 1765308861
transform 1 0 1730 0 1 434
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_3
timestamp 1765308861
transform 1 0 1974 0 1 436
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_4
timestamp 1765308861
transform 1 0 2221 0 1 439
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_5
timestamp 1765308861
transform 1 0 2455 0 1 438
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_6
timestamp 1765308861
transform 1 0 2717 0 1 439
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_7
timestamp 1765308861
transform 1 0 2952 0 1 437
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_8
timestamp 1765308861
transform 1 0 3698 0 1 423
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_9
timestamp 1765308861
transform 1 0 814 0 1 1030
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_10
timestamp 1765308861
transform 1 0 1270 0 1 1026
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_11
timestamp 1765308861
transform 1 0 1486 0 1 1025
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_12
timestamp 1765308861
transform 1 0 1696 0 1 1025
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_13
timestamp 1765308861
transform 1 0 1910 0 1 1028
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_14
timestamp 1765308861
transform 1 0 2136 0 1 1027
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_15
timestamp 1765308861
transform 1 0 2348 0 1 1028
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_16
timestamp 1765308861
transform 1 0 2561 0 1 1031
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_17
timestamp 1765308861
transform 1 0 2778 0 1 1030
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_18
timestamp 1765308861
transform 1 0 3283 0 1 1029
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_19
timestamp 1765308861
transform 1 0 3768 0 1 1025
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_20
timestamp 1765308861
transform 1 0 4799 0 1 1022
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_21
timestamp 1765308861
transform 1 0 5016 0 1 1019
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_22
timestamp 1765308861
transform 1 0 5229 0 1 1017
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_23
timestamp 1765308861
transform 1 0 5437 0 1 1022
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_24
timestamp 1765308861
transform 1 0 5654 0 1 1019
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_25
timestamp 1765308861
transform 1 0 5865 0 1 1022
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_26
timestamp 1765308861
transform 1 0 6083 0 1 1019
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_27
timestamp 1765308861
transform 1 0 6572 0 1 1019
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_28
timestamp 1765308861
transform 1 0 4291 0 1 1020
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_29
timestamp 1765308861
transform 1 0 7063 0 1 1032
box -43 -214 99 -158
use via_cont_2um  via_cont_2um_0
timestamp 1765308861
transform 1 0 696 0 1 -46
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_1
timestamp 1765308861
transform 1 0 1450 0 1 -78
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_2
timestamp 1765308861
transform 1 0 1938 0 1 -82
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_3
timestamp 1765308861
transform 1 0 2423 0 1 -75
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_4
timestamp 1765308861
transform 1 0 2916 0 1 -77
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_5
timestamp 1765308861
transform 1 0 766 0 1 1035
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_6
timestamp 1765308861
transform 1 0 972 0 1 1035
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_7
timestamp 1765308861
transform 1 0 1263 0 1 1035
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_8
timestamp 1765308861
transform 1 0 1698 0 1 1034
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_9
timestamp 1765308861
transform 1 0 2127 0 1 1036
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_10
timestamp 1765308861
transform 1 0 2563 0 1 1041
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_11
timestamp 1765308861
transform 1 0 2987 0 1 1033
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_12
timestamp 1765308861
transform 1 0 3904 0 1 -110
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_13
timestamp 1765308861
transform 1 0 4273 0 1 1029
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_14
timestamp 1765308861
transform 1 0 3493 0 1 1041
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_15
timestamp 1765308861
transform 1 0 3774 0 1 1038
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_16
timestamp 1765308861
transform 1 0 4016 0 1 1044
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_17
timestamp 1765308861
transform 1 0 4780 0 1 1032
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_18
timestamp 1765308861
transform 1 0 5211 0 1 1035
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_19
timestamp 1765308861
transform 1 0 5637 0 1 1035
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_20
timestamp 1765308861
transform 1 0 6064 0 1 1040
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_21
timestamp 1765308861
transform 1 0 7070 0 1 1038
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_22
timestamp 1765308861
transform 1 0 6784 0 1 1058
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_23
timestamp 1765308861
transform 1 0 4499 0 1 1030
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_24
timestamp 1765308861
transform 1 0 7288 0 1 1038
box -92 -99 -36 240
use nmos_6p0_B4TB5U  XM0
timestamp 1765308861
transform 1 0 754 0 1 -4
box -334 -432 334 432
use pmos_6p0_CYEQN4  XM1
timestamp 1765308861
transform 1 0 3815 0 1 1093
box -368 -486 378 486
use pmos_6p0_CYEQN4  XM3
timestamp 1765308861
transform 1 0 806 0 1 1093
box -368 -486 378 486
use pmos_6p0_CYEQN4  XM4
timestamp 1765308861
transform 1 0 3313 0 1 1093
box -368 -486 378 486
use pmos_6p0_CYEQN4  XM7
timestamp 1765308861
transform 1 0 6605 0 1 1093
box -368 -486 378 486
use pmos_6p0_CYEQN4  XM9
timestamp 1765308861
transform 1 0 4317 0 1 1093
box -368 -486 378 486
<< labels >>
flabel metal1 s 412 1527 612 1727 0 FreeSans 1600 0 0 0 VDD
port 1 nsew
flabel metal1 s 404 -608 604 -408 0 FreeSans 1600 0 0 0 VSS
port 2 nsew
flabel metal1 s 7380 273 7580 473 0 FreeSans 1600 0 0 0 Vout
port 3 nsew
<< properties >>
string GDS_END 224696
string GDS_FILE ../gds/simple_por.gds.gz
string GDS_START 187224
<< end >>
