magic
tech gf180mcuD
magscale 1 10
timestamp 1765308861
<< pwell >>
rect -334 -432 334 432
<< hvnmos >>
rect -70 -224 70 176
<< mvndiff >>
rect -158 140 -70 176
rect -158 -188 -145 140
rect -99 -188 -70 140
rect -158 -224 -70 -188
rect 70 140 158 176
rect 70 -188 99 140
rect 145 -188 158 140
rect 70 -224 158 -188
<< mvndiffc >>
rect -145 -188 -99 140
rect 99 -188 145 140
<< mvpsubdiff >>
rect -302 328 302 400
rect -302 258 -230 328
rect -302 -258 -289 258
rect -243 -258 -230 258
rect 230 258 302 328
rect -302 -328 -230 -258
rect 230 -258 243 258
rect 289 -258 302 258
rect 230 -328 302 -258
rect -302 -341 302 -328
rect -302 -387 -164 -341
rect 164 -387 302 -341
rect -302 -400 302 -387
<< mvpsubdiffcont >>
rect -289 -258 -243 258
rect 243 -258 289 258
rect -164 -387 164 -341
<< polysilicon >>
rect -70 255 70 268
rect -70 209 -23 255
rect 23 209 70 255
rect -70 176 70 209
rect -70 -268 70 -224
<< polycontact >>
rect -23 209 23 255
<< metal1 >>
rect -289 341 289 387
rect -289 258 -243 341
rect 243 258 289 341
rect -68 209 -23 255
rect 23 209 68 255
rect -145 140 -99 174
rect -145 -222 -99 -188
rect 99 140 145 174
rect 99 -222 145 -188
rect -289 -341 -243 -258
rect 243 -341 289 -258
rect -289 -387 -164 -341
rect 164 -387 289 -341
<< properties >>
string FIXED_BBOX -266 -364 266 364
string GDS_END 30080
string GDS_FILE ../gds/simple_por.gds.gz
string GDS_START 26684
<< end >>
