magic
tech gf180mcuD
magscale 1 10
timestamp 1765308861
<< metal1 >>
rect 3923 8645 6463 8714
rect 3923 8593 3979 8645
rect 4031 8593 4103 8645
rect 4155 8593 4227 8645
rect 4279 8593 4351 8645
rect 4403 8593 4475 8645
rect 4527 8593 4599 8645
rect 4651 8593 4723 8645
rect 4775 8593 4847 8645
rect 4899 8593 4971 8645
rect 5023 8593 5095 8645
rect 5147 8593 5219 8645
rect 5271 8593 5343 8645
rect 5395 8593 5467 8645
rect 5519 8593 5591 8645
rect 5643 8593 5715 8645
rect 5767 8593 5839 8645
rect 5891 8593 5963 8645
rect 6015 8593 6087 8645
rect 6139 8593 6211 8645
rect 6263 8593 6335 8645
rect 6387 8593 6463 8645
rect 3923 8521 6463 8593
rect 3923 8469 3979 8521
rect 4031 8469 4103 8521
rect 4155 8469 4227 8521
rect 4279 8469 4351 8521
rect 4403 8469 4475 8521
rect 4527 8469 4599 8521
rect 4651 8469 4723 8521
rect 4775 8469 4847 8521
rect 4899 8469 4971 8521
rect 5023 8469 5095 8521
rect 5147 8469 5219 8521
rect 5271 8469 5343 8521
rect 5395 8469 5467 8521
rect 5519 8469 5591 8521
rect 5643 8469 5715 8521
rect 5767 8469 5839 8521
rect 5891 8469 5963 8521
rect 6015 8469 6087 8521
rect 6139 8469 6211 8521
rect 6263 8469 6335 8521
rect 6387 8469 6463 8521
rect 3923 8397 6463 8469
rect 3923 8345 3979 8397
rect 4031 8345 4103 8397
rect 4155 8345 4227 8397
rect 4279 8345 4351 8397
rect 4403 8345 4475 8397
rect 4527 8345 4599 8397
rect 4651 8345 4723 8397
rect 4775 8345 4847 8397
rect 4899 8345 4971 8397
rect 5023 8345 5095 8397
rect 5147 8345 5219 8397
rect 5271 8345 5343 8397
rect 5395 8345 5467 8397
rect 5519 8345 5591 8397
rect 5643 8345 5715 8397
rect 5767 8345 5839 8397
rect 5891 8345 5963 8397
rect 6015 8345 6087 8397
rect 6139 8345 6211 8397
rect 6263 8345 6335 8397
rect 6387 8345 6463 8397
rect 3923 8273 6463 8345
rect 3923 8221 3979 8273
rect 4031 8221 4103 8273
rect 4155 8221 4227 8273
rect 4279 8221 4351 8273
rect 4403 8221 4475 8273
rect 4527 8221 4599 8273
rect 4651 8221 4723 8273
rect 4775 8221 4847 8273
rect 4899 8221 4971 8273
rect 5023 8221 5095 8273
rect 5147 8221 5219 8273
rect 5271 8221 5343 8273
rect 5395 8221 5467 8273
rect 5519 8221 5591 8273
rect 5643 8221 5715 8273
rect 5767 8221 5839 8273
rect 5891 8221 5963 8273
rect 6015 8221 6087 8273
rect 6139 8221 6211 8273
rect 6263 8221 6335 8273
rect 6387 8221 6463 8273
rect 3923 8149 6463 8221
rect 3923 8097 3979 8149
rect 4031 8097 4103 8149
rect 4155 8097 4227 8149
rect 4279 8097 4351 8149
rect 4403 8097 4475 8149
rect 4527 8097 4599 8149
rect 4651 8097 4723 8149
rect 4775 8097 4847 8149
rect 4899 8097 4971 8149
rect 5023 8097 5095 8149
rect 5147 8097 5219 8149
rect 5271 8097 5343 8149
rect 5395 8097 5467 8149
rect 5519 8097 5591 8149
rect 5643 8097 5715 8149
rect 5767 8097 5839 8149
rect 5891 8097 5963 8149
rect 6015 8097 6087 8149
rect 6139 8097 6211 8149
rect 6263 8097 6335 8149
rect 6387 8097 6463 8149
rect 3923 8025 6463 8097
rect 20890 8226 21090 8247
rect 20890 8070 20911 8226
rect 21067 8070 21090 8226
rect 20890 8047 21090 8070
rect 22253 8206 22453 8227
rect 22253 8050 22274 8206
rect 22430 8050 22453 8206
rect 3923 7973 3979 8025
rect 4031 7973 4103 8025
rect 4155 7973 4227 8025
rect 4279 7973 4351 8025
rect 4403 7973 4475 8025
rect 4527 7973 4599 8025
rect 4651 7973 4723 8025
rect 4775 7973 4847 8025
rect 4899 7973 4971 8025
rect 5023 7973 5095 8025
rect 5147 7973 5219 8025
rect 5271 7973 5343 8025
rect 5395 7973 5467 8025
rect 5519 7973 5591 8025
rect 5643 7973 5715 8025
rect 5767 7973 5839 8025
rect 5891 7973 5963 8025
rect 6015 7973 6087 8025
rect 6139 7973 6211 8025
rect 6263 7973 6335 8025
rect 6387 7973 6463 8025
rect 3923 7914 6463 7973
rect 20642 7959 20643 7974
rect 20907 7959 21045 8047
rect 22253 8027 22453 8050
rect 20642 7831 21045 7959
rect 20907 6821 21045 7831
rect 22342 7592 22451 8027
rect 3953 6625 6493 6684
rect 3953 6573 4019 6625
rect 4071 6573 4143 6625
rect 4195 6573 4267 6625
rect 4319 6573 4391 6625
rect 4443 6573 4515 6625
rect 4567 6573 4639 6625
rect 4691 6573 4763 6625
rect 4815 6573 4887 6625
rect 4939 6573 5011 6625
rect 5063 6573 5135 6625
rect 5187 6573 5259 6625
rect 5311 6573 5383 6625
rect 5435 6573 5507 6625
rect 5559 6573 5631 6625
rect 5683 6573 5755 6625
rect 5807 6573 5879 6625
rect 5931 6573 6003 6625
rect 6055 6573 6127 6625
rect 6179 6573 6251 6625
rect 6303 6573 6375 6625
rect 6427 6573 6493 6625
rect 3953 6501 6493 6573
rect 3953 6449 4019 6501
rect 4071 6449 4143 6501
rect 4195 6449 4267 6501
rect 4319 6449 4391 6501
rect 4443 6449 4515 6501
rect 4567 6449 4639 6501
rect 4691 6449 4763 6501
rect 4815 6449 4887 6501
rect 4939 6449 5011 6501
rect 5063 6449 5135 6501
rect 5187 6449 5259 6501
rect 5311 6449 5383 6501
rect 5435 6449 5507 6501
rect 5559 6449 5631 6501
rect 5683 6449 5755 6501
rect 5807 6449 5879 6501
rect 5931 6449 6003 6501
rect 6055 6449 6127 6501
rect 6179 6449 6251 6501
rect 6303 6449 6375 6501
rect 6427 6449 6493 6501
rect 3953 6377 6493 6449
rect 3953 6325 4019 6377
rect 4071 6325 4143 6377
rect 4195 6325 4267 6377
rect 4319 6325 4391 6377
rect 4443 6325 4515 6377
rect 4567 6325 4639 6377
rect 4691 6325 4763 6377
rect 4815 6325 4887 6377
rect 4939 6325 5011 6377
rect 5063 6325 5135 6377
rect 5187 6325 5259 6377
rect 5311 6325 5383 6377
rect 5435 6325 5507 6377
rect 5559 6325 5631 6377
rect 5683 6325 5755 6377
rect 5807 6325 5879 6377
rect 5931 6325 6003 6377
rect 6055 6325 6127 6377
rect 6179 6325 6251 6377
rect 6303 6325 6375 6377
rect 6427 6325 6493 6377
rect 22096 6567 22204 7023
rect 22342 6808 22452 7592
rect 24708 6995 24908 7017
rect 24085 6994 24908 6995
rect 24085 6838 24730 6994
rect 24886 6838 24908 6994
rect 24085 6826 24908 6838
rect 24708 6817 24908 6826
rect 22096 6546 22310 6567
rect 22096 6390 22131 6546
rect 22287 6390 22310 6546
rect 22096 6367 22310 6390
rect 23960 6529 24160 6544
rect 24709 6529 24909 6542
rect 23960 6523 24909 6529
rect 23960 6367 23981 6523
rect 24137 6521 24909 6523
rect 24137 6367 24731 6521
rect 23960 6365 24731 6367
rect 24887 6365 24909 6521
rect 23960 6360 24909 6365
rect 23960 6344 24160 6360
rect 24709 6342 24909 6360
rect 3953 6253 6493 6325
rect 3953 6201 4019 6253
rect 4071 6201 4143 6253
rect 4195 6201 4267 6253
rect 4319 6201 4391 6253
rect 4443 6201 4515 6253
rect 4567 6201 4639 6253
rect 4691 6201 4763 6253
rect 4815 6201 4887 6253
rect 4939 6201 5011 6253
rect 5063 6201 5135 6253
rect 5187 6201 5259 6253
rect 5311 6201 5383 6253
rect 5435 6201 5507 6253
rect 5559 6201 5631 6253
rect 5683 6201 5755 6253
rect 5807 6201 5879 6253
rect 5931 6201 6003 6253
rect 6055 6201 6127 6253
rect 6179 6201 6251 6253
rect 6303 6201 6375 6253
rect 6427 6201 6493 6253
rect 3953 6129 6493 6201
rect 3953 6077 4019 6129
rect 4071 6077 4143 6129
rect 4195 6077 4267 6129
rect 4319 6077 4391 6129
rect 4443 6077 4515 6129
rect 4567 6077 4639 6129
rect 4691 6077 4763 6129
rect 4815 6077 4887 6129
rect 4939 6077 5011 6129
rect 5063 6077 5135 6129
rect 5187 6077 5259 6129
rect 5311 6077 5383 6129
rect 5435 6077 5507 6129
rect 5559 6077 5631 6129
rect 5683 6077 5755 6129
rect 5807 6077 5879 6129
rect 5931 6077 6003 6129
rect 6055 6077 6127 6129
rect 6179 6077 6251 6129
rect 6303 6077 6375 6129
rect 6427 6077 6493 6129
rect 3953 6005 6493 6077
rect 3953 5953 4019 6005
rect 4071 5953 4143 6005
rect 4195 5953 4267 6005
rect 4319 5953 4391 6005
rect 4443 5953 4515 6005
rect 4567 5953 4639 6005
rect 4691 5953 4763 6005
rect 4815 5953 4887 6005
rect 4939 5953 5011 6005
rect 5063 5953 5135 6005
rect 5187 5953 5259 6005
rect 5311 5953 5383 6005
rect 5435 5953 5507 6005
rect 5559 5953 5631 6005
rect 5683 5953 5755 6005
rect 5807 5953 5879 6005
rect 5931 5953 6003 6005
rect 6055 5953 6127 6005
rect 6179 5953 6251 6005
rect 6303 5953 6375 6005
rect 6427 5953 6493 6005
rect 3953 5884 6493 5953
<< via1 >>
rect 3979 8593 4031 8645
rect 4103 8593 4155 8645
rect 4227 8593 4279 8645
rect 4351 8593 4403 8645
rect 4475 8593 4527 8645
rect 4599 8593 4651 8645
rect 4723 8593 4775 8645
rect 4847 8593 4899 8645
rect 4971 8593 5023 8645
rect 5095 8593 5147 8645
rect 5219 8593 5271 8645
rect 5343 8593 5395 8645
rect 5467 8593 5519 8645
rect 5591 8593 5643 8645
rect 5715 8593 5767 8645
rect 5839 8593 5891 8645
rect 5963 8593 6015 8645
rect 6087 8593 6139 8645
rect 6211 8593 6263 8645
rect 6335 8593 6387 8645
rect 3979 8469 4031 8521
rect 4103 8469 4155 8521
rect 4227 8469 4279 8521
rect 4351 8469 4403 8521
rect 4475 8469 4527 8521
rect 4599 8469 4651 8521
rect 4723 8469 4775 8521
rect 4847 8469 4899 8521
rect 4971 8469 5023 8521
rect 5095 8469 5147 8521
rect 5219 8469 5271 8521
rect 5343 8469 5395 8521
rect 5467 8469 5519 8521
rect 5591 8469 5643 8521
rect 5715 8469 5767 8521
rect 5839 8469 5891 8521
rect 5963 8469 6015 8521
rect 6087 8469 6139 8521
rect 6211 8469 6263 8521
rect 6335 8469 6387 8521
rect 3979 8345 4031 8397
rect 4103 8345 4155 8397
rect 4227 8345 4279 8397
rect 4351 8345 4403 8397
rect 4475 8345 4527 8397
rect 4599 8345 4651 8397
rect 4723 8345 4775 8397
rect 4847 8345 4899 8397
rect 4971 8345 5023 8397
rect 5095 8345 5147 8397
rect 5219 8345 5271 8397
rect 5343 8345 5395 8397
rect 5467 8345 5519 8397
rect 5591 8345 5643 8397
rect 5715 8345 5767 8397
rect 5839 8345 5891 8397
rect 5963 8345 6015 8397
rect 6087 8345 6139 8397
rect 6211 8345 6263 8397
rect 6335 8345 6387 8397
rect 3979 8221 4031 8273
rect 4103 8221 4155 8273
rect 4227 8221 4279 8273
rect 4351 8221 4403 8273
rect 4475 8221 4527 8273
rect 4599 8221 4651 8273
rect 4723 8221 4775 8273
rect 4847 8221 4899 8273
rect 4971 8221 5023 8273
rect 5095 8221 5147 8273
rect 5219 8221 5271 8273
rect 5343 8221 5395 8273
rect 5467 8221 5519 8273
rect 5591 8221 5643 8273
rect 5715 8221 5767 8273
rect 5839 8221 5891 8273
rect 5963 8221 6015 8273
rect 6087 8221 6139 8273
rect 6211 8221 6263 8273
rect 6335 8221 6387 8273
rect 3979 8097 4031 8149
rect 4103 8097 4155 8149
rect 4227 8097 4279 8149
rect 4351 8097 4403 8149
rect 4475 8097 4527 8149
rect 4599 8097 4651 8149
rect 4723 8097 4775 8149
rect 4847 8097 4899 8149
rect 4971 8097 5023 8149
rect 5095 8097 5147 8149
rect 5219 8097 5271 8149
rect 5343 8097 5395 8149
rect 5467 8097 5519 8149
rect 5591 8097 5643 8149
rect 5715 8097 5767 8149
rect 5839 8097 5891 8149
rect 5963 8097 6015 8149
rect 6087 8097 6139 8149
rect 6211 8097 6263 8149
rect 6335 8097 6387 8149
rect 20911 8070 21067 8226
rect 22274 8050 22430 8206
rect 3979 7973 4031 8025
rect 4103 7973 4155 8025
rect 4227 7973 4279 8025
rect 4351 7973 4403 8025
rect 4475 7973 4527 8025
rect 4599 7973 4651 8025
rect 4723 7973 4775 8025
rect 4847 7973 4899 8025
rect 4971 7973 5023 8025
rect 5095 7973 5147 8025
rect 5219 7973 5271 8025
rect 5343 7973 5395 8025
rect 5467 7973 5519 8025
rect 5591 7973 5643 8025
rect 5715 7973 5767 8025
rect 5839 7973 5891 8025
rect 5963 7973 6015 8025
rect 6087 7973 6139 8025
rect 6211 7973 6263 8025
rect 6335 7973 6387 8025
rect 4019 6573 4071 6625
rect 4143 6573 4195 6625
rect 4267 6573 4319 6625
rect 4391 6573 4443 6625
rect 4515 6573 4567 6625
rect 4639 6573 4691 6625
rect 4763 6573 4815 6625
rect 4887 6573 4939 6625
rect 5011 6573 5063 6625
rect 5135 6573 5187 6625
rect 5259 6573 5311 6625
rect 5383 6573 5435 6625
rect 5507 6573 5559 6625
rect 5631 6573 5683 6625
rect 5755 6573 5807 6625
rect 5879 6573 5931 6625
rect 6003 6573 6055 6625
rect 6127 6573 6179 6625
rect 6251 6573 6303 6625
rect 6375 6573 6427 6625
rect 4019 6449 4071 6501
rect 4143 6449 4195 6501
rect 4267 6449 4319 6501
rect 4391 6449 4443 6501
rect 4515 6449 4567 6501
rect 4639 6449 4691 6501
rect 4763 6449 4815 6501
rect 4887 6449 4939 6501
rect 5011 6449 5063 6501
rect 5135 6449 5187 6501
rect 5259 6449 5311 6501
rect 5383 6449 5435 6501
rect 5507 6449 5559 6501
rect 5631 6449 5683 6501
rect 5755 6449 5807 6501
rect 5879 6449 5931 6501
rect 6003 6449 6055 6501
rect 6127 6449 6179 6501
rect 6251 6449 6303 6501
rect 6375 6449 6427 6501
rect 4019 6325 4071 6377
rect 4143 6325 4195 6377
rect 4267 6325 4319 6377
rect 4391 6325 4443 6377
rect 4515 6325 4567 6377
rect 4639 6325 4691 6377
rect 4763 6325 4815 6377
rect 4887 6325 4939 6377
rect 5011 6325 5063 6377
rect 5135 6325 5187 6377
rect 5259 6325 5311 6377
rect 5383 6325 5435 6377
rect 5507 6325 5559 6377
rect 5631 6325 5683 6377
rect 5755 6325 5807 6377
rect 5879 6325 5931 6377
rect 6003 6325 6055 6377
rect 6127 6325 6179 6377
rect 6251 6325 6303 6377
rect 6375 6325 6427 6377
rect 24730 6838 24886 6994
rect 22131 6390 22287 6546
rect 23981 6367 24137 6523
rect 24731 6365 24887 6521
rect 4019 6201 4071 6253
rect 4143 6201 4195 6253
rect 4267 6201 4319 6253
rect 4391 6201 4443 6253
rect 4515 6201 4567 6253
rect 4639 6201 4691 6253
rect 4763 6201 4815 6253
rect 4887 6201 4939 6253
rect 5011 6201 5063 6253
rect 5135 6201 5187 6253
rect 5259 6201 5311 6253
rect 5383 6201 5435 6253
rect 5507 6201 5559 6253
rect 5631 6201 5683 6253
rect 5755 6201 5807 6253
rect 5879 6201 5931 6253
rect 6003 6201 6055 6253
rect 6127 6201 6179 6253
rect 6251 6201 6303 6253
rect 6375 6201 6427 6253
rect 4019 6077 4071 6129
rect 4143 6077 4195 6129
rect 4267 6077 4319 6129
rect 4391 6077 4443 6129
rect 4515 6077 4567 6129
rect 4639 6077 4691 6129
rect 4763 6077 4815 6129
rect 4887 6077 4939 6129
rect 5011 6077 5063 6129
rect 5135 6077 5187 6129
rect 5259 6077 5311 6129
rect 5383 6077 5435 6129
rect 5507 6077 5559 6129
rect 5631 6077 5683 6129
rect 5755 6077 5807 6129
rect 5879 6077 5931 6129
rect 6003 6077 6055 6129
rect 6127 6077 6179 6129
rect 6251 6077 6303 6129
rect 6375 6077 6427 6129
rect 4019 5953 4071 6005
rect 4143 5953 4195 6005
rect 4267 5953 4319 6005
rect 4391 5953 4443 6005
rect 4515 5953 4567 6005
rect 4639 5953 4691 6005
rect 4763 5953 4815 6005
rect 4887 5953 4939 6005
rect 5011 5953 5063 6005
rect 5135 5953 5187 6005
rect 5259 5953 5311 6005
rect 5383 5953 5435 6005
rect 5507 5953 5559 6005
rect 5631 5953 5683 6005
rect 5755 5953 5807 6005
rect 5879 5953 5931 6005
rect 6003 5953 6055 6005
rect 6127 5953 6179 6005
rect 6251 5953 6303 6005
rect 6375 5953 6427 6005
<< metal2 >>
rect 3923 8647 6463 8714
rect 3923 8591 3977 8647
rect 4033 8591 4101 8647
rect 4157 8591 4225 8647
rect 4281 8591 4349 8647
rect 4405 8591 4473 8647
rect 4529 8591 4597 8647
rect 4653 8591 4721 8647
rect 4777 8591 4845 8647
rect 4901 8591 4969 8647
rect 5025 8591 5093 8647
rect 5149 8591 5217 8647
rect 5273 8591 5341 8647
rect 5397 8591 5465 8647
rect 5521 8591 5589 8647
rect 5645 8591 5713 8647
rect 5769 8591 5837 8647
rect 5893 8591 5961 8647
rect 6017 8591 6085 8647
rect 6141 8591 6209 8647
rect 6265 8591 6333 8647
rect 6389 8591 6463 8647
rect 3923 8523 6463 8591
rect 3923 8467 3977 8523
rect 4033 8467 4101 8523
rect 4157 8467 4225 8523
rect 4281 8467 4349 8523
rect 4405 8467 4473 8523
rect 4529 8467 4597 8523
rect 4653 8467 4721 8523
rect 4777 8467 4845 8523
rect 4901 8467 4969 8523
rect 5025 8467 5093 8523
rect 5149 8467 5217 8523
rect 5273 8467 5341 8523
rect 5397 8467 5465 8523
rect 5521 8467 5589 8523
rect 5645 8467 5713 8523
rect 5769 8467 5837 8523
rect 5893 8467 5961 8523
rect 6017 8467 6085 8523
rect 6141 8467 6209 8523
rect 6265 8467 6333 8523
rect 6389 8467 6463 8523
rect 3923 8399 6463 8467
rect 3923 8343 3977 8399
rect 4033 8343 4101 8399
rect 4157 8343 4225 8399
rect 4281 8343 4349 8399
rect 4405 8343 4473 8399
rect 4529 8343 4597 8399
rect 4653 8343 4721 8399
rect 4777 8343 4845 8399
rect 4901 8343 4969 8399
rect 5025 8343 5093 8399
rect 5149 8343 5217 8399
rect 5273 8343 5341 8399
rect 5397 8343 5465 8399
rect 5521 8343 5589 8399
rect 5645 8343 5713 8399
rect 5769 8343 5837 8399
rect 5893 8343 5961 8399
rect 6017 8343 6085 8399
rect 6141 8343 6209 8399
rect 6265 8343 6333 8399
rect 6389 8343 6463 8399
rect 3923 8275 6463 8343
rect 3923 8219 3977 8275
rect 4033 8219 4101 8275
rect 4157 8219 4225 8275
rect 4281 8219 4349 8275
rect 4405 8219 4473 8275
rect 4529 8219 4597 8275
rect 4653 8219 4721 8275
rect 4777 8219 4845 8275
rect 4901 8219 4969 8275
rect 5025 8219 5093 8275
rect 5149 8219 5217 8275
rect 5273 8219 5341 8275
rect 5397 8219 5465 8275
rect 5521 8219 5589 8275
rect 5645 8219 5713 8275
rect 5769 8219 5837 8275
rect 5893 8219 5961 8275
rect 6017 8219 6085 8275
rect 6141 8219 6209 8275
rect 6265 8219 6333 8275
rect 6389 8219 6463 8275
rect 20948 8465 22404 8602
rect 20948 8247 21085 8465
rect 3923 8151 6463 8219
rect 3923 8095 3977 8151
rect 4033 8095 4101 8151
rect 4157 8095 4225 8151
rect 4281 8095 4349 8151
rect 4405 8095 4473 8151
rect 4529 8095 4597 8151
rect 4653 8095 4721 8151
rect 4777 8095 4845 8151
rect 4901 8095 4969 8151
rect 5025 8095 5093 8151
rect 5149 8095 5217 8151
rect 5273 8095 5341 8151
rect 5397 8095 5465 8151
rect 5521 8095 5589 8151
rect 5645 8095 5713 8151
rect 5769 8095 5837 8151
rect 5893 8095 5961 8151
rect 6017 8095 6085 8151
rect 6141 8095 6209 8151
rect 6265 8095 6333 8151
rect 6389 8095 6463 8151
rect 3923 8027 6463 8095
rect 20890 8226 21090 8247
rect 22267 8227 22404 8465
rect 20890 8070 20911 8226
rect 21067 8070 21090 8226
rect 20890 8047 21090 8070
rect 22253 8206 22453 8227
rect 22253 8050 22274 8206
rect 22430 8050 22453 8206
rect 22253 8027 22453 8050
rect 3923 7971 3977 8027
rect 4033 7971 4101 8027
rect 4157 7971 4225 8027
rect 4281 7971 4349 8027
rect 4405 7971 4473 8027
rect 4529 7971 4597 8027
rect 4653 7971 4721 8027
rect 4777 7971 4845 8027
rect 4901 7971 4969 8027
rect 5025 7971 5093 8027
rect 5149 7971 5217 8027
rect 5273 7971 5341 8027
rect 5397 7971 5465 8027
rect 5521 7971 5589 8027
rect 5645 7971 5713 8027
rect 5769 7971 5837 8027
rect 5893 7971 5961 8027
rect 6017 7971 6085 8027
rect 6141 7971 6209 8027
rect 6265 7971 6333 8027
rect 6389 7971 6463 8027
rect 3923 7914 6463 7971
rect 7152 7602 7520 7647
rect 3953 6627 6493 6684
rect 3953 6571 4017 6627
rect 4073 6571 4141 6627
rect 4197 6571 4265 6627
rect 4321 6571 4389 6627
rect 4445 6571 4513 6627
rect 4569 6571 4637 6627
rect 4693 6571 4761 6627
rect 4817 6571 4885 6627
rect 4941 6571 5009 6627
rect 5065 6571 5133 6627
rect 5189 6571 5257 6627
rect 5313 6571 5381 6627
rect 5437 6571 5505 6627
rect 5561 6571 5629 6627
rect 5685 6571 5753 6627
rect 5809 6571 5877 6627
rect 5933 6571 6001 6627
rect 6057 6571 6125 6627
rect 6181 6571 6249 6627
rect 6305 6571 6373 6627
rect 6429 6571 6493 6627
rect 3953 6503 6493 6571
rect 7152 6610 7199 7602
rect 7463 6610 7520 7602
rect 7152 6561 7520 6610
rect 17284 7458 17907 7555
rect 17284 7402 17377 7458
rect 17433 7402 17501 7458
rect 17557 7402 17625 7458
rect 17681 7402 17749 7458
rect 17805 7402 17907 7458
rect 17284 7334 17907 7402
rect 17284 7278 17377 7334
rect 17433 7278 17501 7334
rect 17557 7278 17625 7334
rect 17681 7278 17749 7334
rect 17805 7278 17907 7334
rect 17284 7210 17907 7278
rect 17284 7154 17377 7210
rect 17433 7154 17501 7210
rect 17557 7154 17625 7210
rect 17681 7154 17749 7210
rect 17805 7154 17907 7210
rect 17284 7086 17907 7154
rect 17284 7030 17377 7086
rect 17433 7030 17501 7086
rect 17557 7030 17625 7086
rect 17681 7030 17749 7086
rect 17805 7030 17907 7086
rect 17284 6962 17907 7030
rect 17284 6906 17377 6962
rect 17433 6906 17501 6962
rect 17557 6906 17625 6962
rect 17681 6906 17749 6962
rect 17805 6906 17907 6962
rect 17284 6857 17907 6906
rect 24708 6994 25108 7017
rect 17284 6838 18224 6857
rect 17284 6782 17377 6838
rect 17433 6782 17501 6838
rect 17557 6782 17625 6838
rect 17681 6782 17749 6838
rect 17805 6782 18224 6838
rect 24708 6838 24730 6994
rect 24886 6838 25108 6994
rect 24708 6817 25108 6838
rect 17284 6714 18224 6782
rect 17284 6658 17377 6714
rect 17433 6658 17501 6714
rect 17557 6658 17625 6714
rect 17681 6658 17749 6714
rect 17805 6659 18224 6714
rect 17805 6658 17907 6659
rect 17284 6590 17907 6658
rect 3953 6447 4017 6503
rect 4073 6447 4141 6503
rect 4197 6447 4265 6503
rect 4321 6447 4389 6503
rect 4445 6447 4513 6503
rect 4569 6447 4637 6503
rect 4693 6447 4761 6503
rect 4817 6447 4885 6503
rect 4941 6447 5009 6503
rect 5065 6447 5133 6503
rect 5189 6447 5257 6503
rect 5313 6447 5381 6503
rect 5437 6447 5505 6503
rect 5561 6447 5629 6503
rect 5685 6447 5753 6503
rect 5809 6447 5877 6503
rect 5933 6447 6001 6503
rect 6057 6447 6125 6503
rect 6181 6447 6249 6503
rect 6305 6447 6373 6503
rect 6429 6447 6493 6503
rect 3953 6379 6493 6447
rect 3953 6323 4017 6379
rect 4073 6323 4141 6379
rect 4197 6323 4265 6379
rect 4321 6323 4389 6379
rect 4445 6323 4513 6379
rect 4569 6323 4637 6379
rect 4693 6323 4761 6379
rect 4817 6323 4885 6379
rect 4941 6323 5009 6379
rect 5065 6323 5133 6379
rect 5189 6323 5257 6379
rect 5313 6323 5381 6379
rect 5437 6323 5505 6379
rect 5561 6323 5629 6379
rect 5685 6323 5753 6379
rect 5809 6323 5877 6379
rect 5933 6323 6001 6379
rect 6057 6323 6125 6379
rect 6181 6323 6249 6379
rect 6305 6323 6373 6379
rect 6429 6323 6493 6379
rect 3953 6255 6493 6323
rect 17284 6534 17377 6590
rect 17433 6534 17501 6590
rect 17557 6534 17625 6590
rect 17681 6534 17749 6590
rect 17805 6534 17907 6590
rect 17284 6466 17907 6534
rect 17284 6410 17377 6466
rect 17433 6410 17501 6466
rect 17557 6410 17625 6466
rect 17681 6410 17749 6466
rect 17805 6410 17907 6466
rect 17284 6306 17907 6410
rect 22110 6546 22310 6567
rect 22110 6390 22131 6546
rect 22287 6390 22310 6546
rect 22110 6367 22310 6390
rect 23960 6523 24160 6544
rect 23960 6367 23981 6523
rect 24137 6367 24160 6523
rect 3953 6199 4017 6255
rect 4073 6199 4141 6255
rect 4197 6199 4265 6255
rect 4321 6199 4389 6255
rect 4445 6199 4513 6255
rect 4569 6199 4637 6255
rect 4693 6199 4761 6255
rect 4817 6199 4885 6255
rect 4941 6199 5009 6255
rect 5065 6199 5133 6255
rect 5189 6199 5257 6255
rect 5313 6199 5381 6255
rect 5437 6199 5505 6255
rect 5561 6199 5629 6255
rect 5685 6199 5753 6255
rect 5809 6199 5877 6255
rect 5933 6199 6001 6255
rect 6057 6199 6125 6255
rect 6181 6199 6249 6255
rect 6305 6199 6373 6255
rect 6429 6199 6493 6255
rect 3953 6131 6493 6199
rect 3953 6075 4017 6131
rect 4073 6075 4141 6131
rect 4197 6075 4265 6131
rect 4321 6075 4389 6131
rect 4445 6075 4513 6131
rect 4569 6075 4637 6131
rect 4693 6075 4761 6131
rect 4817 6075 4885 6131
rect 4941 6075 5009 6131
rect 5065 6075 5133 6131
rect 5189 6075 5257 6131
rect 5313 6075 5381 6131
rect 5437 6075 5505 6131
rect 5561 6075 5629 6131
rect 5685 6075 5753 6131
rect 5809 6075 5877 6131
rect 5933 6075 6001 6131
rect 6057 6075 6125 6131
rect 6181 6075 6249 6131
rect 6305 6075 6373 6131
rect 6429 6075 6493 6131
rect 3953 6007 6493 6075
rect 3953 5951 4017 6007
rect 4073 5951 4141 6007
rect 4197 5951 4265 6007
rect 4321 5951 4389 6007
rect 4445 5951 4513 6007
rect 4569 5951 4637 6007
rect 4693 5951 4761 6007
rect 4817 5951 4885 6007
rect 4941 5951 5009 6007
rect 5065 5951 5133 6007
rect 5189 5951 5257 6007
rect 5313 5951 5381 6007
rect 5437 5951 5505 6007
rect 5561 5951 5629 6007
rect 5685 5951 5753 6007
rect 5809 5951 5877 6007
rect 5933 5951 6001 6007
rect 6057 5951 6125 6007
rect 6181 5951 6249 6007
rect 6305 5951 6373 6007
rect 6429 5951 6493 6007
rect 3953 5884 6493 5951
rect 22185 5910 22306 6367
rect 23960 6344 24160 6367
rect 24709 6521 25109 6542
rect 24709 6365 24731 6521
rect 24887 6365 25109 6521
rect 23989 5910 24125 6344
rect 24709 6342 25109 6365
rect 22185 5774 24125 5910
<< via2 >>
rect 3977 8645 4033 8647
rect 3977 8593 3979 8645
rect 3979 8593 4031 8645
rect 4031 8593 4033 8645
rect 3977 8591 4033 8593
rect 4101 8645 4157 8647
rect 4101 8593 4103 8645
rect 4103 8593 4155 8645
rect 4155 8593 4157 8645
rect 4101 8591 4157 8593
rect 4225 8645 4281 8647
rect 4225 8593 4227 8645
rect 4227 8593 4279 8645
rect 4279 8593 4281 8645
rect 4225 8591 4281 8593
rect 4349 8645 4405 8647
rect 4349 8593 4351 8645
rect 4351 8593 4403 8645
rect 4403 8593 4405 8645
rect 4349 8591 4405 8593
rect 4473 8645 4529 8647
rect 4473 8593 4475 8645
rect 4475 8593 4527 8645
rect 4527 8593 4529 8645
rect 4473 8591 4529 8593
rect 4597 8645 4653 8647
rect 4597 8593 4599 8645
rect 4599 8593 4651 8645
rect 4651 8593 4653 8645
rect 4597 8591 4653 8593
rect 4721 8645 4777 8647
rect 4721 8593 4723 8645
rect 4723 8593 4775 8645
rect 4775 8593 4777 8645
rect 4721 8591 4777 8593
rect 4845 8645 4901 8647
rect 4845 8593 4847 8645
rect 4847 8593 4899 8645
rect 4899 8593 4901 8645
rect 4845 8591 4901 8593
rect 4969 8645 5025 8647
rect 4969 8593 4971 8645
rect 4971 8593 5023 8645
rect 5023 8593 5025 8645
rect 4969 8591 5025 8593
rect 5093 8645 5149 8647
rect 5093 8593 5095 8645
rect 5095 8593 5147 8645
rect 5147 8593 5149 8645
rect 5093 8591 5149 8593
rect 5217 8645 5273 8647
rect 5217 8593 5219 8645
rect 5219 8593 5271 8645
rect 5271 8593 5273 8645
rect 5217 8591 5273 8593
rect 5341 8645 5397 8647
rect 5341 8593 5343 8645
rect 5343 8593 5395 8645
rect 5395 8593 5397 8645
rect 5341 8591 5397 8593
rect 5465 8645 5521 8647
rect 5465 8593 5467 8645
rect 5467 8593 5519 8645
rect 5519 8593 5521 8645
rect 5465 8591 5521 8593
rect 5589 8645 5645 8647
rect 5589 8593 5591 8645
rect 5591 8593 5643 8645
rect 5643 8593 5645 8645
rect 5589 8591 5645 8593
rect 5713 8645 5769 8647
rect 5713 8593 5715 8645
rect 5715 8593 5767 8645
rect 5767 8593 5769 8645
rect 5713 8591 5769 8593
rect 5837 8645 5893 8647
rect 5837 8593 5839 8645
rect 5839 8593 5891 8645
rect 5891 8593 5893 8645
rect 5837 8591 5893 8593
rect 5961 8645 6017 8647
rect 5961 8593 5963 8645
rect 5963 8593 6015 8645
rect 6015 8593 6017 8645
rect 5961 8591 6017 8593
rect 6085 8645 6141 8647
rect 6085 8593 6087 8645
rect 6087 8593 6139 8645
rect 6139 8593 6141 8645
rect 6085 8591 6141 8593
rect 6209 8645 6265 8647
rect 6209 8593 6211 8645
rect 6211 8593 6263 8645
rect 6263 8593 6265 8645
rect 6209 8591 6265 8593
rect 6333 8645 6389 8647
rect 6333 8593 6335 8645
rect 6335 8593 6387 8645
rect 6387 8593 6389 8645
rect 6333 8591 6389 8593
rect 3977 8521 4033 8523
rect 3977 8469 3979 8521
rect 3979 8469 4031 8521
rect 4031 8469 4033 8521
rect 3977 8467 4033 8469
rect 4101 8521 4157 8523
rect 4101 8469 4103 8521
rect 4103 8469 4155 8521
rect 4155 8469 4157 8521
rect 4101 8467 4157 8469
rect 4225 8521 4281 8523
rect 4225 8469 4227 8521
rect 4227 8469 4279 8521
rect 4279 8469 4281 8521
rect 4225 8467 4281 8469
rect 4349 8521 4405 8523
rect 4349 8469 4351 8521
rect 4351 8469 4403 8521
rect 4403 8469 4405 8521
rect 4349 8467 4405 8469
rect 4473 8521 4529 8523
rect 4473 8469 4475 8521
rect 4475 8469 4527 8521
rect 4527 8469 4529 8521
rect 4473 8467 4529 8469
rect 4597 8521 4653 8523
rect 4597 8469 4599 8521
rect 4599 8469 4651 8521
rect 4651 8469 4653 8521
rect 4597 8467 4653 8469
rect 4721 8521 4777 8523
rect 4721 8469 4723 8521
rect 4723 8469 4775 8521
rect 4775 8469 4777 8521
rect 4721 8467 4777 8469
rect 4845 8521 4901 8523
rect 4845 8469 4847 8521
rect 4847 8469 4899 8521
rect 4899 8469 4901 8521
rect 4845 8467 4901 8469
rect 4969 8521 5025 8523
rect 4969 8469 4971 8521
rect 4971 8469 5023 8521
rect 5023 8469 5025 8521
rect 4969 8467 5025 8469
rect 5093 8521 5149 8523
rect 5093 8469 5095 8521
rect 5095 8469 5147 8521
rect 5147 8469 5149 8521
rect 5093 8467 5149 8469
rect 5217 8521 5273 8523
rect 5217 8469 5219 8521
rect 5219 8469 5271 8521
rect 5271 8469 5273 8521
rect 5217 8467 5273 8469
rect 5341 8521 5397 8523
rect 5341 8469 5343 8521
rect 5343 8469 5395 8521
rect 5395 8469 5397 8521
rect 5341 8467 5397 8469
rect 5465 8521 5521 8523
rect 5465 8469 5467 8521
rect 5467 8469 5519 8521
rect 5519 8469 5521 8521
rect 5465 8467 5521 8469
rect 5589 8521 5645 8523
rect 5589 8469 5591 8521
rect 5591 8469 5643 8521
rect 5643 8469 5645 8521
rect 5589 8467 5645 8469
rect 5713 8521 5769 8523
rect 5713 8469 5715 8521
rect 5715 8469 5767 8521
rect 5767 8469 5769 8521
rect 5713 8467 5769 8469
rect 5837 8521 5893 8523
rect 5837 8469 5839 8521
rect 5839 8469 5891 8521
rect 5891 8469 5893 8521
rect 5837 8467 5893 8469
rect 5961 8521 6017 8523
rect 5961 8469 5963 8521
rect 5963 8469 6015 8521
rect 6015 8469 6017 8521
rect 5961 8467 6017 8469
rect 6085 8521 6141 8523
rect 6085 8469 6087 8521
rect 6087 8469 6139 8521
rect 6139 8469 6141 8521
rect 6085 8467 6141 8469
rect 6209 8521 6265 8523
rect 6209 8469 6211 8521
rect 6211 8469 6263 8521
rect 6263 8469 6265 8521
rect 6209 8467 6265 8469
rect 6333 8521 6389 8523
rect 6333 8469 6335 8521
rect 6335 8469 6387 8521
rect 6387 8469 6389 8521
rect 6333 8467 6389 8469
rect 3977 8397 4033 8399
rect 3977 8345 3979 8397
rect 3979 8345 4031 8397
rect 4031 8345 4033 8397
rect 3977 8343 4033 8345
rect 4101 8397 4157 8399
rect 4101 8345 4103 8397
rect 4103 8345 4155 8397
rect 4155 8345 4157 8397
rect 4101 8343 4157 8345
rect 4225 8397 4281 8399
rect 4225 8345 4227 8397
rect 4227 8345 4279 8397
rect 4279 8345 4281 8397
rect 4225 8343 4281 8345
rect 4349 8397 4405 8399
rect 4349 8345 4351 8397
rect 4351 8345 4403 8397
rect 4403 8345 4405 8397
rect 4349 8343 4405 8345
rect 4473 8397 4529 8399
rect 4473 8345 4475 8397
rect 4475 8345 4527 8397
rect 4527 8345 4529 8397
rect 4473 8343 4529 8345
rect 4597 8397 4653 8399
rect 4597 8345 4599 8397
rect 4599 8345 4651 8397
rect 4651 8345 4653 8397
rect 4597 8343 4653 8345
rect 4721 8397 4777 8399
rect 4721 8345 4723 8397
rect 4723 8345 4775 8397
rect 4775 8345 4777 8397
rect 4721 8343 4777 8345
rect 4845 8397 4901 8399
rect 4845 8345 4847 8397
rect 4847 8345 4899 8397
rect 4899 8345 4901 8397
rect 4845 8343 4901 8345
rect 4969 8397 5025 8399
rect 4969 8345 4971 8397
rect 4971 8345 5023 8397
rect 5023 8345 5025 8397
rect 4969 8343 5025 8345
rect 5093 8397 5149 8399
rect 5093 8345 5095 8397
rect 5095 8345 5147 8397
rect 5147 8345 5149 8397
rect 5093 8343 5149 8345
rect 5217 8397 5273 8399
rect 5217 8345 5219 8397
rect 5219 8345 5271 8397
rect 5271 8345 5273 8397
rect 5217 8343 5273 8345
rect 5341 8397 5397 8399
rect 5341 8345 5343 8397
rect 5343 8345 5395 8397
rect 5395 8345 5397 8397
rect 5341 8343 5397 8345
rect 5465 8397 5521 8399
rect 5465 8345 5467 8397
rect 5467 8345 5519 8397
rect 5519 8345 5521 8397
rect 5465 8343 5521 8345
rect 5589 8397 5645 8399
rect 5589 8345 5591 8397
rect 5591 8345 5643 8397
rect 5643 8345 5645 8397
rect 5589 8343 5645 8345
rect 5713 8397 5769 8399
rect 5713 8345 5715 8397
rect 5715 8345 5767 8397
rect 5767 8345 5769 8397
rect 5713 8343 5769 8345
rect 5837 8397 5893 8399
rect 5837 8345 5839 8397
rect 5839 8345 5891 8397
rect 5891 8345 5893 8397
rect 5837 8343 5893 8345
rect 5961 8397 6017 8399
rect 5961 8345 5963 8397
rect 5963 8345 6015 8397
rect 6015 8345 6017 8397
rect 5961 8343 6017 8345
rect 6085 8397 6141 8399
rect 6085 8345 6087 8397
rect 6087 8345 6139 8397
rect 6139 8345 6141 8397
rect 6085 8343 6141 8345
rect 6209 8397 6265 8399
rect 6209 8345 6211 8397
rect 6211 8345 6263 8397
rect 6263 8345 6265 8397
rect 6209 8343 6265 8345
rect 6333 8397 6389 8399
rect 6333 8345 6335 8397
rect 6335 8345 6387 8397
rect 6387 8345 6389 8397
rect 6333 8343 6389 8345
rect 3977 8273 4033 8275
rect 3977 8221 3979 8273
rect 3979 8221 4031 8273
rect 4031 8221 4033 8273
rect 3977 8219 4033 8221
rect 4101 8273 4157 8275
rect 4101 8221 4103 8273
rect 4103 8221 4155 8273
rect 4155 8221 4157 8273
rect 4101 8219 4157 8221
rect 4225 8273 4281 8275
rect 4225 8221 4227 8273
rect 4227 8221 4279 8273
rect 4279 8221 4281 8273
rect 4225 8219 4281 8221
rect 4349 8273 4405 8275
rect 4349 8221 4351 8273
rect 4351 8221 4403 8273
rect 4403 8221 4405 8273
rect 4349 8219 4405 8221
rect 4473 8273 4529 8275
rect 4473 8221 4475 8273
rect 4475 8221 4527 8273
rect 4527 8221 4529 8273
rect 4473 8219 4529 8221
rect 4597 8273 4653 8275
rect 4597 8221 4599 8273
rect 4599 8221 4651 8273
rect 4651 8221 4653 8273
rect 4597 8219 4653 8221
rect 4721 8273 4777 8275
rect 4721 8221 4723 8273
rect 4723 8221 4775 8273
rect 4775 8221 4777 8273
rect 4721 8219 4777 8221
rect 4845 8273 4901 8275
rect 4845 8221 4847 8273
rect 4847 8221 4899 8273
rect 4899 8221 4901 8273
rect 4845 8219 4901 8221
rect 4969 8273 5025 8275
rect 4969 8221 4971 8273
rect 4971 8221 5023 8273
rect 5023 8221 5025 8273
rect 4969 8219 5025 8221
rect 5093 8273 5149 8275
rect 5093 8221 5095 8273
rect 5095 8221 5147 8273
rect 5147 8221 5149 8273
rect 5093 8219 5149 8221
rect 5217 8273 5273 8275
rect 5217 8221 5219 8273
rect 5219 8221 5271 8273
rect 5271 8221 5273 8273
rect 5217 8219 5273 8221
rect 5341 8273 5397 8275
rect 5341 8221 5343 8273
rect 5343 8221 5395 8273
rect 5395 8221 5397 8273
rect 5341 8219 5397 8221
rect 5465 8273 5521 8275
rect 5465 8221 5467 8273
rect 5467 8221 5519 8273
rect 5519 8221 5521 8273
rect 5465 8219 5521 8221
rect 5589 8273 5645 8275
rect 5589 8221 5591 8273
rect 5591 8221 5643 8273
rect 5643 8221 5645 8273
rect 5589 8219 5645 8221
rect 5713 8273 5769 8275
rect 5713 8221 5715 8273
rect 5715 8221 5767 8273
rect 5767 8221 5769 8273
rect 5713 8219 5769 8221
rect 5837 8273 5893 8275
rect 5837 8221 5839 8273
rect 5839 8221 5891 8273
rect 5891 8221 5893 8273
rect 5837 8219 5893 8221
rect 5961 8273 6017 8275
rect 5961 8221 5963 8273
rect 5963 8221 6015 8273
rect 6015 8221 6017 8273
rect 5961 8219 6017 8221
rect 6085 8273 6141 8275
rect 6085 8221 6087 8273
rect 6087 8221 6139 8273
rect 6139 8221 6141 8273
rect 6085 8219 6141 8221
rect 6209 8273 6265 8275
rect 6209 8221 6211 8273
rect 6211 8221 6263 8273
rect 6263 8221 6265 8273
rect 6209 8219 6265 8221
rect 6333 8273 6389 8275
rect 6333 8221 6335 8273
rect 6335 8221 6387 8273
rect 6387 8221 6389 8273
rect 6333 8219 6389 8221
rect 3977 8149 4033 8151
rect 3977 8097 3979 8149
rect 3979 8097 4031 8149
rect 4031 8097 4033 8149
rect 3977 8095 4033 8097
rect 4101 8149 4157 8151
rect 4101 8097 4103 8149
rect 4103 8097 4155 8149
rect 4155 8097 4157 8149
rect 4101 8095 4157 8097
rect 4225 8149 4281 8151
rect 4225 8097 4227 8149
rect 4227 8097 4279 8149
rect 4279 8097 4281 8149
rect 4225 8095 4281 8097
rect 4349 8149 4405 8151
rect 4349 8097 4351 8149
rect 4351 8097 4403 8149
rect 4403 8097 4405 8149
rect 4349 8095 4405 8097
rect 4473 8149 4529 8151
rect 4473 8097 4475 8149
rect 4475 8097 4527 8149
rect 4527 8097 4529 8149
rect 4473 8095 4529 8097
rect 4597 8149 4653 8151
rect 4597 8097 4599 8149
rect 4599 8097 4651 8149
rect 4651 8097 4653 8149
rect 4597 8095 4653 8097
rect 4721 8149 4777 8151
rect 4721 8097 4723 8149
rect 4723 8097 4775 8149
rect 4775 8097 4777 8149
rect 4721 8095 4777 8097
rect 4845 8149 4901 8151
rect 4845 8097 4847 8149
rect 4847 8097 4899 8149
rect 4899 8097 4901 8149
rect 4845 8095 4901 8097
rect 4969 8149 5025 8151
rect 4969 8097 4971 8149
rect 4971 8097 5023 8149
rect 5023 8097 5025 8149
rect 4969 8095 5025 8097
rect 5093 8149 5149 8151
rect 5093 8097 5095 8149
rect 5095 8097 5147 8149
rect 5147 8097 5149 8149
rect 5093 8095 5149 8097
rect 5217 8149 5273 8151
rect 5217 8097 5219 8149
rect 5219 8097 5271 8149
rect 5271 8097 5273 8149
rect 5217 8095 5273 8097
rect 5341 8149 5397 8151
rect 5341 8097 5343 8149
rect 5343 8097 5395 8149
rect 5395 8097 5397 8149
rect 5341 8095 5397 8097
rect 5465 8149 5521 8151
rect 5465 8097 5467 8149
rect 5467 8097 5519 8149
rect 5519 8097 5521 8149
rect 5465 8095 5521 8097
rect 5589 8149 5645 8151
rect 5589 8097 5591 8149
rect 5591 8097 5643 8149
rect 5643 8097 5645 8149
rect 5589 8095 5645 8097
rect 5713 8149 5769 8151
rect 5713 8097 5715 8149
rect 5715 8097 5767 8149
rect 5767 8097 5769 8149
rect 5713 8095 5769 8097
rect 5837 8149 5893 8151
rect 5837 8097 5839 8149
rect 5839 8097 5891 8149
rect 5891 8097 5893 8149
rect 5837 8095 5893 8097
rect 5961 8149 6017 8151
rect 5961 8097 5963 8149
rect 5963 8097 6015 8149
rect 6015 8097 6017 8149
rect 5961 8095 6017 8097
rect 6085 8149 6141 8151
rect 6085 8097 6087 8149
rect 6087 8097 6139 8149
rect 6139 8097 6141 8149
rect 6085 8095 6141 8097
rect 6209 8149 6265 8151
rect 6209 8097 6211 8149
rect 6211 8097 6263 8149
rect 6263 8097 6265 8149
rect 6209 8095 6265 8097
rect 6333 8149 6389 8151
rect 6333 8097 6335 8149
rect 6335 8097 6387 8149
rect 6387 8097 6389 8149
rect 6333 8095 6389 8097
rect 3977 8025 4033 8027
rect 3977 7973 3979 8025
rect 3979 7973 4031 8025
rect 4031 7973 4033 8025
rect 3977 7971 4033 7973
rect 4101 8025 4157 8027
rect 4101 7973 4103 8025
rect 4103 7973 4155 8025
rect 4155 7973 4157 8025
rect 4101 7971 4157 7973
rect 4225 8025 4281 8027
rect 4225 7973 4227 8025
rect 4227 7973 4279 8025
rect 4279 7973 4281 8025
rect 4225 7971 4281 7973
rect 4349 8025 4405 8027
rect 4349 7973 4351 8025
rect 4351 7973 4403 8025
rect 4403 7973 4405 8025
rect 4349 7971 4405 7973
rect 4473 8025 4529 8027
rect 4473 7973 4475 8025
rect 4475 7973 4527 8025
rect 4527 7973 4529 8025
rect 4473 7971 4529 7973
rect 4597 8025 4653 8027
rect 4597 7973 4599 8025
rect 4599 7973 4651 8025
rect 4651 7973 4653 8025
rect 4597 7971 4653 7973
rect 4721 8025 4777 8027
rect 4721 7973 4723 8025
rect 4723 7973 4775 8025
rect 4775 7973 4777 8025
rect 4721 7971 4777 7973
rect 4845 8025 4901 8027
rect 4845 7973 4847 8025
rect 4847 7973 4899 8025
rect 4899 7973 4901 8025
rect 4845 7971 4901 7973
rect 4969 8025 5025 8027
rect 4969 7973 4971 8025
rect 4971 7973 5023 8025
rect 5023 7973 5025 8025
rect 4969 7971 5025 7973
rect 5093 8025 5149 8027
rect 5093 7973 5095 8025
rect 5095 7973 5147 8025
rect 5147 7973 5149 8025
rect 5093 7971 5149 7973
rect 5217 8025 5273 8027
rect 5217 7973 5219 8025
rect 5219 7973 5271 8025
rect 5271 7973 5273 8025
rect 5217 7971 5273 7973
rect 5341 8025 5397 8027
rect 5341 7973 5343 8025
rect 5343 7973 5395 8025
rect 5395 7973 5397 8025
rect 5341 7971 5397 7973
rect 5465 8025 5521 8027
rect 5465 7973 5467 8025
rect 5467 7973 5519 8025
rect 5519 7973 5521 8025
rect 5465 7971 5521 7973
rect 5589 8025 5645 8027
rect 5589 7973 5591 8025
rect 5591 7973 5643 8025
rect 5643 7973 5645 8025
rect 5589 7971 5645 7973
rect 5713 8025 5769 8027
rect 5713 7973 5715 8025
rect 5715 7973 5767 8025
rect 5767 7973 5769 8025
rect 5713 7971 5769 7973
rect 5837 8025 5893 8027
rect 5837 7973 5839 8025
rect 5839 7973 5891 8025
rect 5891 7973 5893 8025
rect 5837 7971 5893 7973
rect 5961 8025 6017 8027
rect 5961 7973 5963 8025
rect 5963 7973 6015 8025
rect 6015 7973 6017 8025
rect 5961 7971 6017 7973
rect 6085 8025 6141 8027
rect 6085 7973 6087 8025
rect 6087 7973 6139 8025
rect 6139 7973 6141 8025
rect 6085 7971 6141 7973
rect 6209 8025 6265 8027
rect 6209 7973 6211 8025
rect 6211 7973 6263 8025
rect 6263 7973 6265 8025
rect 6209 7971 6265 7973
rect 6333 8025 6389 8027
rect 6333 7973 6335 8025
rect 6335 7973 6387 8025
rect 6387 7973 6389 8025
rect 6333 7971 6389 7973
rect 4017 6625 4073 6627
rect 4017 6573 4019 6625
rect 4019 6573 4071 6625
rect 4071 6573 4073 6625
rect 4017 6571 4073 6573
rect 4141 6625 4197 6627
rect 4141 6573 4143 6625
rect 4143 6573 4195 6625
rect 4195 6573 4197 6625
rect 4141 6571 4197 6573
rect 4265 6625 4321 6627
rect 4265 6573 4267 6625
rect 4267 6573 4319 6625
rect 4319 6573 4321 6625
rect 4265 6571 4321 6573
rect 4389 6625 4445 6627
rect 4389 6573 4391 6625
rect 4391 6573 4443 6625
rect 4443 6573 4445 6625
rect 4389 6571 4445 6573
rect 4513 6625 4569 6627
rect 4513 6573 4515 6625
rect 4515 6573 4567 6625
rect 4567 6573 4569 6625
rect 4513 6571 4569 6573
rect 4637 6625 4693 6627
rect 4637 6573 4639 6625
rect 4639 6573 4691 6625
rect 4691 6573 4693 6625
rect 4637 6571 4693 6573
rect 4761 6625 4817 6627
rect 4761 6573 4763 6625
rect 4763 6573 4815 6625
rect 4815 6573 4817 6625
rect 4761 6571 4817 6573
rect 4885 6625 4941 6627
rect 4885 6573 4887 6625
rect 4887 6573 4939 6625
rect 4939 6573 4941 6625
rect 4885 6571 4941 6573
rect 5009 6625 5065 6627
rect 5009 6573 5011 6625
rect 5011 6573 5063 6625
rect 5063 6573 5065 6625
rect 5009 6571 5065 6573
rect 5133 6625 5189 6627
rect 5133 6573 5135 6625
rect 5135 6573 5187 6625
rect 5187 6573 5189 6625
rect 5133 6571 5189 6573
rect 5257 6625 5313 6627
rect 5257 6573 5259 6625
rect 5259 6573 5311 6625
rect 5311 6573 5313 6625
rect 5257 6571 5313 6573
rect 5381 6625 5437 6627
rect 5381 6573 5383 6625
rect 5383 6573 5435 6625
rect 5435 6573 5437 6625
rect 5381 6571 5437 6573
rect 5505 6625 5561 6627
rect 5505 6573 5507 6625
rect 5507 6573 5559 6625
rect 5559 6573 5561 6625
rect 5505 6571 5561 6573
rect 5629 6625 5685 6627
rect 5629 6573 5631 6625
rect 5631 6573 5683 6625
rect 5683 6573 5685 6625
rect 5629 6571 5685 6573
rect 5753 6625 5809 6627
rect 5753 6573 5755 6625
rect 5755 6573 5807 6625
rect 5807 6573 5809 6625
rect 5753 6571 5809 6573
rect 5877 6625 5933 6627
rect 5877 6573 5879 6625
rect 5879 6573 5931 6625
rect 5931 6573 5933 6625
rect 5877 6571 5933 6573
rect 6001 6625 6057 6627
rect 6001 6573 6003 6625
rect 6003 6573 6055 6625
rect 6055 6573 6057 6625
rect 6001 6571 6057 6573
rect 6125 6625 6181 6627
rect 6125 6573 6127 6625
rect 6127 6573 6179 6625
rect 6179 6573 6181 6625
rect 6125 6571 6181 6573
rect 6249 6625 6305 6627
rect 6249 6573 6251 6625
rect 6251 6573 6303 6625
rect 6303 6573 6305 6625
rect 6249 6571 6305 6573
rect 6373 6625 6429 6627
rect 6373 6573 6375 6625
rect 6375 6573 6427 6625
rect 6427 6573 6429 6625
rect 6373 6571 6429 6573
rect 7199 6610 7463 7602
rect 17377 7402 17433 7458
rect 17501 7402 17557 7458
rect 17625 7402 17681 7458
rect 17749 7402 17805 7458
rect 17377 7278 17433 7334
rect 17501 7278 17557 7334
rect 17625 7278 17681 7334
rect 17749 7278 17805 7334
rect 17377 7154 17433 7210
rect 17501 7154 17557 7210
rect 17625 7154 17681 7210
rect 17749 7154 17805 7210
rect 17377 7030 17433 7086
rect 17501 7030 17557 7086
rect 17625 7030 17681 7086
rect 17749 7030 17805 7086
rect 17377 6906 17433 6962
rect 17501 6906 17557 6962
rect 17625 6906 17681 6962
rect 17749 6906 17805 6962
rect 17377 6782 17433 6838
rect 17501 6782 17557 6838
rect 17625 6782 17681 6838
rect 17749 6782 17805 6838
rect 17377 6658 17433 6714
rect 17501 6658 17557 6714
rect 17625 6658 17681 6714
rect 17749 6658 17805 6714
rect 4017 6501 4073 6503
rect 4017 6449 4019 6501
rect 4019 6449 4071 6501
rect 4071 6449 4073 6501
rect 4017 6447 4073 6449
rect 4141 6501 4197 6503
rect 4141 6449 4143 6501
rect 4143 6449 4195 6501
rect 4195 6449 4197 6501
rect 4141 6447 4197 6449
rect 4265 6501 4321 6503
rect 4265 6449 4267 6501
rect 4267 6449 4319 6501
rect 4319 6449 4321 6501
rect 4265 6447 4321 6449
rect 4389 6501 4445 6503
rect 4389 6449 4391 6501
rect 4391 6449 4443 6501
rect 4443 6449 4445 6501
rect 4389 6447 4445 6449
rect 4513 6501 4569 6503
rect 4513 6449 4515 6501
rect 4515 6449 4567 6501
rect 4567 6449 4569 6501
rect 4513 6447 4569 6449
rect 4637 6501 4693 6503
rect 4637 6449 4639 6501
rect 4639 6449 4691 6501
rect 4691 6449 4693 6501
rect 4637 6447 4693 6449
rect 4761 6501 4817 6503
rect 4761 6449 4763 6501
rect 4763 6449 4815 6501
rect 4815 6449 4817 6501
rect 4761 6447 4817 6449
rect 4885 6501 4941 6503
rect 4885 6449 4887 6501
rect 4887 6449 4939 6501
rect 4939 6449 4941 6501
rect 4885 6447 4941 6449
rect 5009 6501 5065 6503
rect 5009 6449 5011 6501
rect 5011 6449 5063 6501
rect 5063 6449 5065 6501
rect 5009 6447 5065 6449
rect 5133 6501 5189 6503
rect 5133 6449 5135 6501
rect 5135 6449 5187 6501
rect 5187 6449 5189 6501
rect 5133 6447 5189 6449
rect 5257 6501 5313 6503
rect 5257 6449 5259 6501
rect 5259 6449 5311 6501
rect 5311 6449 5313 6501
rect 5257 6447 5313 6449
rect 5381 6501 5437 6503
rect 5381 6449 5383 6501
rect 5383 6449 5435 6501
rect 5435 6449 5437 6501
rect 5381 6447 5437 6449
rect 5505 6501 5561 6503
rect 5505 6449 5507 6501
rect 5507 6449 5559 6501
rect 5559 6449 5561 6501
rect 5505 6447 5561 6449
rect 5629 6501 5685 6503
rect 5629 6449 5631 6501
rect 5631 6449 5683 6501
rect 5683 6449 5685 6501
rect 5629 6447 5685 6449
rect 5753 6501 5809 6503
rect 5753 6449 5755 6501
rect 5755 6449 5807 6501
rect 5807 6449 5809 6501
rect 5753 6447 5809 6449
rect 5877 6501 5933 6503
rect 5877 6449 5879 6501
rect 5879 6449 5931 6501
rect 5931 6449 5933 6501
rect 5877 6447 5933 6449
rect 6001 6501 6057 6503
rect 6001 6449 6003 6501
rect 6003 6449 6055 6501
rect 6055 6449 6057 6501
rect 6001 6447 6057 6449
rect 6125 6501 6181 6503
rect 6125 6449 6127 6501
rect 6127 6449 6179 6501
rect 6179 6449 6181 6501
rect 6125 6447 6181 6449
rect 6249 6501 6305 6503
rect 6249 6449 6251 6501
rect 6251 6449 6303 6501
rect 6303 6449 6305 6501
rect 6249 6447 6305 6449
rect 6373 6501 6429 6503
rect 6373 6449 6375 6501
rect 6375 6449 6427 6501
rect 6427 6449 6429 6501
rect 6373 6447 6429 6449
rect 4017 6377 4073 6379
rect 4017 6325 4019 6377
rect 4019 6325 4071 6377
rect 4071 6325 4073 6377
rect 4017 6323 4073 6325
rect 4141 6377 4197 6379
rect 4141 6325 4143 6377
rect 4143 6325 4195 6377
rect 4195 6325 4197 6377
rect 4141 6323 4197 6325
rect 4265 6377 4321 6379
rect 4265 6325 4267 6377
rect 4267 6325 4319 6377
rect 4319 6325 4321 6377
rect 4265 6323 4321 6325
rect 4389 6377 4445 6379
rect 4389 6325 4391 6377
rect 4391 6325 4443 6377
rect 4443 6325 4445 6377
rect 4389 6323 4445 6325
rect 4513 6377 4569 6379
rect 4513 6325 4515 6377
rect 4515 6325 4567 6377
rect 4567 6325 4569 6377
rect 4513 6323 4569 6325
rect 4637 6377 4693 6379
rect 4637 6325 4639 6377
rect 4639 6325 4691 6377
rect 4691 6325 4693 6377
rect 4637 6323 4693 6325
rect 4761 6377 4817 6379
rect 4761 6325 4763 6377
rect 4763 6325 4815 6377
rect 4815 6325 4817 6377
rect 4761 6323 4817 6325
rect 4885 6377 4941 6379
rect 4885 6325 4887 6377
rect 4887 6325 4939 6377
rect 4939 6325 4941 6377
rect 4885 6323 4941 6325
rect 5009 6377 5065 6379
rect 5009 6325 5011 6377
rect 5011 6325 5063 6377
rect 5063 6325 5065 6377
rect 5009 6323 5065 6325
rect 5133 6377 5189 6379
rect 5133 6325 5135 6377
rect 5135 6325 5187 6377
rect 5187 6325 5189 6377
rect 5133 6323 5189 6325
rect 5257 6377 5313 6379
rect 5257 6325 5259 6377
rect 5259 6325 5311 6377
rect 5311 6325 5313 6377
rect 5257 6323 5313 6325
rect 5381 6377 5437 6379
rect 5381 6325 5383 6377
rect 5383 6325 5435 6377
rect 5435 6325 5437 6377
rect 5381 6323 5437 6325
rect 5505 6377 5561 6379
rect 5505 6325 5507 6377
rect 5507 6325 5559 6377
rect 5559 6325 5561 6377
rect 5505 6323 5561 6325
rect 5629 6377 5685 6379
rect 5629 6325 5631 6377
rect 5631 6325 5683 6377
rect 5683 6325 5685 6377
rect 5629 6323 5685 6325
rect 5753 6377 5809 6379
rect 5753 6325 5755 6377
rect 5755 6325 5807 6377
rect 5807 6325 5809 6377
rect 5753 6323 5809 6325
rect 5877 6377 5933 6379
rect 5877 6325 5879 6377
rect 5879 6325 5931 6377
rect 5931 6325 5933 6377
rect 5877 6323 5933 6325
rect 6001 6377 6057 6379
rect 6001 6325 6003 6377
rect 6003 6325 6055 6377
rect 6055 6325 6057 6377
rect 6001 6323 6057 6325
rect 6125 6377 6181 6379
rect 6125 6325 6127 6377
rect 6127 6325 6179 6377
rect 6179 6325 6181 6377
rect 6125 6323 6181 6325
rect 6249 6377 6305 6379
rect 6249 6325 6251 6377
rect 6251 6325 6303 6377
rect 6303 6325 6305 6377
rect 6249 6323 6305 6325
rect 6373 6377 6429 6379
rect 6373 6325 6375 6377
rect 6375 6325 6427 6377
rect 6427 6325 6429 6377
rect 6373 6323 6429 6325
rect 17377 6534 17433 6590
rect 17501 6534 17557 6590
rect 17625 6534 17681 6590
rect 17749 6534 17805 6590
rect 17377 6410 17433 6466
rect 17501 6410 17557 6466
rect 17625 6410 17681 6466
rect 17749 6410 17805 6466
rect 4017 6253 4073 6255
rect 4017 6201 4019 6253
rect 4019 6201 4071 6253
rect 4071 6201 4073 6253
rect 4017 6199 4073 6201
rect 4141 6253 4197 6255
rect 4141 6201 4143 6253
rect 4143 6201 4195 6253
rect 4195 6201 4197 6253
rect 4141 6199 4197 6201
rect 4265 6253 4321 6255
rect 4265 6201 4267 6253
rect 4267 6201 4319 6253
rect 4319 6201 4321 6253
rect 4265 6199 4321 6201
rect 4389 6253 4445 6255
rect 4389 6201 4391 6253
rect 4391 6201 4443 6253
rect 4443 6201 4445 6253
rect 4389 6199 4445 6201
rect 4513 6253 4569 6255
rect 4513 6201 4515 6253
rect 4515 6201 4567 6253
rect 4567 6201 4569 6253
rect 4513 6199 4569 6201
rect 4637 6253 4693 6255
rect 4637 6201 4639 6253
rect 4639 6201 4691 6253
rect 4691 6201 4693 6253
rect 4637 6199 4693 6201
rect 4761 6253 4817 6255
rect 4761 6201 4763 6253
rect 4763 6201 4815 6253
rect 4815 6201 4817 6253
rect 4761 6199 4817 6201
rect 4885 6253 4941 6255
rect 4885 6201 4887 6253
rect 4887 6201 4939 6253
rect 4939 6201 4941 6253
rect 4885 6199 4941 6201
rect 5009 6253 5065 6255
rect 5009 6201 5011 6253
rect 5011 6201 5063 6253
rect 5063 6201 5065 6253
rect 5009 6199 5065 6201
rect 5133 6253 5189 6255
rect 5133 6201 5135 6253
rect 5135 6201 5187 6253
rect 5187 6201 5189 6253
rect 5133 6199 5189 6201
rect 5257 6253 5313 6255
rect 5257 6201 5259 6253
rect 5259 6201 5311 6253
rect 5311 6201 5313 6253
rect 5257 6199 5313 6201
rect 5381 6253 5437 6255
rect 5381 6201 5383 6253
rect 5383 6201 5435 6253
rect 5435 6201 5437 6253
rect 5381 6199 5437 6201
rect 5505 6253 5561 6255
rect 5505 6201 5507 6253
rect 5507 6201 5559 6253
rect 5559 6201 5561 6253
rect 5505 6199 5561 6201
rect 5629 6253 5685 6255
rect 5629 6201 5631 6253
rect 5631 6201 5683 6253
rect 5683 6201 5685 6253
rect 5629 6199 5685 6201
rect 5753 6253 5809 6255
rect 5753 6201 5755 6253
rect 5755 6201 5807 6253
rect 5807 6201 5809 6253
rect 5753 6199 5809 6201
rect 5877 6253 5933 6255
rect 5877 6201 5879 6253
rect 5879 6201 5931 6253
rect 5931 6201 5933 6253
rect 5877 6199 5933 6201
rect 6001 6253 6057 6255
rect 6001 6201 6003 6253
rect 6003 6201 6055 6253
rect 6055 6201 6057 6253
rect 6001 6199 6057 6201
rect 6125 6253 6181 6255
rect 6125 6201 6127 6253
rect 6127 6201 6179 6253
rect 6179 6201 6181 6253
rect 6125 6199 6181 6201
rect 6249 6253 6305 6255
rect 6249 6201 6251 6253
rect 6251 6201 6303 6253
rect 6303 6201 6305 6253
rect 6249 6199 6305 6201
rect 6373 6253 6429 6255
rect 6373 6201 6375 6253
rect 6375 6201 6427 6253
rect 6427 6201 6429 6253
rect 6373 6199 6429 6201
rect 4017 6129 4073 6131
rect 4017 6077 4019 6129
rect 4019 6077 4071 6129
rect 4071 6077 4073 6129
rect 4017 6075 4073 6077
rect 4141 6129 4197 6131
rect 4141 6077 4143 6129
rect 4143 6077 4195 6129
rect 4195 6077 4197 6129
rect 4141 6075 4197 6077
rect 4265 6129 4321 6131
rect 4265 6077 4267 6129
rect 4267 6077 4319 6129
rect 4319 6077 4321 6129
rect 4265 6075 4321 6077
rect 4389 6129 4445 6131
rect 4389 6077 4391 6129
rect 4391 6077 4443 6129
rect 4443 6077 4445 6129
rect 4389 6075 4445 6077
rect 4513 6129 4569 6131
rect 4513 6077 4515 6129
rect 4515 6077 4567 6129
rect 4567 6077 4569 6129
rect 4513 6075 4569 6077
rect 4637 6129 4693 6131
rect 4637 6077 4639 6129
rect 4639 6077 4691 6129
rect 4691 6077 4693 6129
rect 4637 6075 4693 6077
rect 4761 6129 4817 6131
rect 4761 6077 4763 6129
rect 4763 6077 4815 6129
rect 4815 6077 4817 6129
rect 4761 6075 4817 6077
rect 4885 6129 4941 6131
rect 4885 6077 4887 6129
rect 4887 6077 4939 6129
rect 4939 6077 4941 6129
rect 4885 6075 4941 6077
rect 5009 6129 5065 6131
rect 5009 6077 5011 6129
rect 5011 6077 5063 6129
rect 5063 6077 5065 6129
rect 5009 6075 5065 6077
rect 5133 6129 5189 6131
rect 5133 6077 5135 6129
rect 5135 6077 5187 6129
rect 5187 6077 5189 6129
rect 5133 6075 5189 6077
rect 5257 6129 5313 6131
rect 5257 6077 5259 6129
rect 5259 6077 5311 6129
rect 5311 6077 5313 6129
rect 5257 6075 5313 6077
rect 5381 6129 5437 6131
rect 5381 6077 5383 6129
rect 5383 6077 5435 6129
rect 5435 6077 5437 6129
rect 5381 6075 5437 6077
rect 5505 6129 5561 6131
rect 5505 6077 5507 6129
rect 5507 6077 5559 6129
rect 5559 6077 5561 6129
rect 5505 6075 5561 6077
rect 5629 6129 5685 6131
rect 5629 6077 5631 6129
rect 5631 6077 5683 6129
rect 5683 6077 5685 6129
rect 5629 6075 5685 6077
rect 5753 6129 5809 6131
rect 5753 6077 5755 6129
rect 5755 6077 5807 6129
rect 5807 6077 5809 6129
rect 5753 6075 5809 6077
rect 5877 6129 5933 6131
rect 5877 6077 5879 6129
rect 5879 6077 5931 6129
rect 5931 6077 5933 6129
rect 5877 6075 5933 6077
rect 6001 6129 6057 6131
rect 6001 6077 6003 6129
rect 6003 6077 6055 6129
rect 6055 6077 6057 6129
rect 6001 6075 6057 6077
rect 6125 6129 6181 6131
rect 6125 6077 6127 6129
rect 6127 6077 6179 6129
rect 6179 6077 6181 6129
rect 6125 6075 6181 6077
rect 6249 6129 6305 6131
rect 6249 6077 6251 6129
rect 6251 6077 6303 6129
rect 6303 6077 6305 6129
rect 6249 6075 6305 6077
rect 6373 6129 6429 6131
rect 6373 6077 6375 6129
rect 6375 6077 6427 6129
rect 6427 6077 6429 6129
rect 6373 6075 6429 6077
rect 4017 6005 4073 6007
rect 4017 5953 4019 6005
rect 4019 5953 4071 6005
rect 4071 5953 4073 6005
rect 4017 5951 4073 5953
rect 4141 6005 4197 6007
rect 4141 5953 4143 6005
rect 4143 5953 4195 6005
rect 4195 5953 4197 6005
rect 4141 5951 4197 5953
rect 4265 6005 4321 6007
rect 4265 5953 4267 6005
rect 4267 5953 4319 6005
rect 4319 5953 4321 6005
rect 4265 5951 4321 5953
rect 4389 6005 4445 6007
rect 4389 5953 4391 6005
rect 4391 5953 4443 6005
rect 4443 5953 4445 6005
rect 4389 5951 4445 5953
rect 4513 6005 4569 6007
rect 4513 5953 4515 6005
rect 4515 5953 4567 6005
rect 4567 5953 4569 6005
rect 4513 5951 4569 5953
rect 4637 6005 4693 6007
rect 4637 5953 4639 6005
rect 4639 5953 4691 6005
rect 4691 5953 4693 6005
rect 4637 5951 4693 5953
rect 4761 6005 4817 6007
rect 4761 5953 4763 6005
rect 4763 5953 4815 6005
rect 4815 5953 4817 6005
rect 4761 5951 4817 5953
rect 4885 6005 4941 6007
rect 4885 5953 4887 6005
rect 4887 5953 4939 6005
rect 4939 5953 4941 6005
rect 4885 5951 4941 5953
rect 5009 6005 5065 6007
rect 5009 5953 5011 6005
rect 5011 5953 5063 6005
rect 5063 5953 5065 6005
rect 5009 5951 5065 5953
rect 5133 6005 5189 6007
rect 5133 5953 5135 6005
rect 5135 5953 5187 6005
rect 5187 5953 5189 6005
rect 5133 5951 5189 5953
rect 5257 6005 5313 6007
rect 5257 5953 5259 6005
rect 5259 5953 5311 6005
rect 5311 5953 5313 6005
rect 5257 5951 5313 5953
rect 5381 6005 5437 6007
rect 5381 5953 5383 6005
rect 5383 5953 5435 6005
rect 5435 5953 5437 6005
rect 5381 5951 5437 5953
rect 5505 6005 5561 6007
rect 5505 5953 5507 6005
rect 5507 5953 5559 6005
rect 5559 5953 5561 6005
rect 5505 5951 5561 5953
rect 5629 6005 5685 6007
rect 5629 5953 5631 6005
rect 5631 5953 5683 6005
rect 5683 5953 5685 6005
rect 5629 5951 5685 5953
rect 5753 6005 5809 6007
rect 5753 5953 5755 6005
rect 5755 5953 5807 6005
rect 5807 5953 5809 6005
rect 5753 5951 5809 5953
rect 5877 6005 5933 6007
rect 5877 5953 5879 6005
rect 5879 5953 5931 6005
rect 5931 5953 5933 6005
rect 5877 5951 5933 5953
rect 6001 6005 6057 6007
rect 6001 5953 6003 6005
rect 6003 5953 6055 6005
rect 6055 5953 6057 6005
rect 6001 5951 6057 5953
rect 6125 6005 6181 6007
rect 6125 5953 6127 6005
rect 6127 5953 6179 6005
rect 6179 5953 6181 6005
rect 6125 5951 6181 5953
rect 6249 6005 6305 6007
rect 6249 5953 6251 6005
rect 6251 5953 6303 6005
rect 6303 5953 6305 6005
rect 6249 5951 6305 5953
rect 6373 6005 6429 6007
rect 6373 5953 6375 6005
rect 6375 5953 6427 6005
rect 6427 5953 6429 6005
rect 6373 5951 6429 5953
<< metal3 >>
rect 3923 8647 6463 8714
rect 3923 8591 3977 8647
rect 4033 8591 4101 8647
rect 4157 8591 4225 8647
rect 4281 8591 4349 8647
rect 4405 8591 4473 8647
rect 4529 8591 4597 8647
rect 4653 8591 4721 8647
rect 4777 8591 4845 8647
rect 4901 8591 4969 8647
rect 5025 8591 5093 8647
rect 5149 8591 5217 8647
rect 5273 8591 5341 8647
rect 5397 8591 5465 8647
rect 5521 8591 5589 8647
rect 5645 8591 5713 8647
rect 5769 8591 5837 8647
rect 5893 8591 5961 8647
rect 6017 8591 6085 8647
rect 6141 8591 6209 8647
rect 6265 8591 6333 8647
rect 6389 8591 6463 8647
rect 3923 8523 6463 8591
rect 3923 8467 3977 8523
rect 4033 8467 4101 8523
rect 4157 8467 4225 8523
rect 4281 8467 4349 8523
rect 4405 8467 4473 8523
rect 4529 8467 4597 8523
rect 4653 8467 4721 8523
rect 4777 8467 4845 8523
rect 4901 8467 4969 8523
rect 5025 8467 5093 8523
rect 5149 8467 5217 8523
rect 5273 8467 5341 8523
rect 5397 8467 5465 8523
rect 5521 8467 5589 8523
rect 5645 8467 5713 8523
rect 5769 8467 5837 8523
rect 5893 8467 5961 8523
rect 6017 8467 6085 8523
rect 6141 8467 6209 8523
rect 6265 8467 6333 8523
rect 6389 8467 6463 8523
rect 3923 8399 6463 8467
rect 3923 8343 3977 8399
rect 4033 8343 4101 8399
rect 4157 8343 4225 8399
rect 4281 8343 4349 8399
rect 4405 8343 4473 8399
rect 4529 8343 4597 8399
rect 4653 8343 4721 8399
rect 4777 8343 4845 8399
rect 4901 8343 4969 8399
rect 5025 8343 5093 8399
rect 5149 8343 5217 8399
rect 5273 8343 5341 8399
rect 5397 8343 5465 8399
rect 5521 8343 5589 8399
rect 5645 8343 5713 8399
rect 5769 8343 5837 8399
rect 5893 8343 5961 8399
rect 6017 8343 6085 8399
rect 6141 8343 6209 8399
rect 6265 8343 6333 8399
rect 6389 8343 6463 8399
rect 3923 8275 6463 8343
rect 3923 8219 3977 8275
rect 4033 8219 4101 8275
rect 4157 8219 4225 8275
rect 4281 8219 4349 8275
rect 4405 8219 4473 8275
rect 4529 8219 4597 8275
rect 4653 8219 4721 8275
rect 4777 8219 4845 8275
rect 4901 8219 4969 8275
rect 5025 8219 5093 8275
rect 5149 8219 5217 8275
rect 5273 8219 5341 8275
rect 5397 8219 5465 8275
rect 5521 8219 5589 8275
rect 5645 8219 5713 8275
rect 5769 8219 5837 8275
rect 5893 8219 5961 8275
rect 6017 8219 6085 8275
rect 6141 8219 6209 8275
rect 6265 8219 6333 8275
rect 6389 8219 6463 8275
rect 3923 8151 6463 8219
rect 3923 8095 3977 8151
rect 4033 8095 4101 8151
rect 4157 8095 4225 8151
rect 4281 8095 4349 8151
rect 4405 8095 4473 8151
rect 4529 8095 4597 8151
rect 4653 8095 4721 8151
rect 4777 8095 4845 8151
rect 4901 8095 4969 8151
rect 5025 8095 5093 8151
rect 5149 8095 5217 8151
rect 5273 8095 5341 8151
rect 5397 8095 5465 8151
rect 5521 8095 5589 8151
rect 5645 8095 5713 8151
rect 5769 8095 5837 8151
rect 5893 8095 5961 8151
rect 6017 8095 6085 8151
rect 6141 8095 6209 8151
rect 6265 8095 6333 8151
rect 6389 8095 6463 8151
rect 3923 8027 6463 8095
rect 3923 7971 3977 8027
rect 4033 7971 4101 8027
rect 4157 7971 4225 8027
rect 4281 7971 4349 8027
rect 4405 7971 4473 8027
rect 4529 7971 4597 8027
rect 4653 7971 4721 8027
rect 4777 7971 4845 8027
rect 4901 7971 4969 8027
rect 5025 7971 5093 8027
rect 5149 7971 5217 8027
rect 5273 7971 5341 8027
rect 5397 7971 5465 8027
rect 5521 7971 5589 8027
rect 5645 7971 5713 8027
rect 5769 7971 5837 8027
rect 5893 7971 5961 8027
rect 6017 7971 6085 8027
rect 6141 7971 6209 8027
rect 6265 7971 6333 8027
rect 6389 7971 6463 8027
rect 3923 7914 6463 7971
rect 7045 7602 7520 7647
rect 3953 6627 6493 6684
rect 3953 6571 4017 6627
rect 4073 6571 4141 6627
rect 4197 6571 4265 6627
rect 4321 6571 4389 6627
rect 4445 6571 4513 6627
rect 4569 6571 4637 6627
rect 4693 6571 4761 6627
rect 4817 6571 4885 6627
rect 4941 6571 5009 6627
rect 5065 6571 5133 6627
rect 5189 6571 5257 6627
rect 5313 6571 5381 6627
rect 5437 6571 5505 6627
rect 5561 6571 5629 6627
rect 5685 6571 5753 6627
rect 5809 6571 5877 6627
rect 5933 6571 6001 6627
rect 6057 6571 6125 6627
rect 6181 6571 6249 6627
rect 6305 6571 6373 6627
rect 6429 6571 6493 6627
rect 3953 6503 6493 6571
rect 7045 6610 7093 7602
rect 7463 6610 7520 7602
rect 7045 6561 7520 6610
rect 17284 7458 17907 7555
rect 17284 7402 17377 7458
rect 17433 7402 17501 7458
rect 17557 7402 17625 7458
rect 17681 7402 17749 7458
rect 17805 7402 17907 7458
rect 17284 7334 17907 7402
rect 17284 7278 17377 7334
rect 17433 7278 17501 7334
rect 17557 7278 17625 7334
rect 17681 7278 17749 7334
rect 17805 7278 17907 7334
rect 17284 7210 17907 7278
rect 17284 7154 17377 7210
rect 17433 7154 17501 7210
rect 17557 7154 17625 7210
rect 17681 7154 17749 7210
rect 17805 7154 17907 7210
rect 17284 7086 17907 7154
rect 17284 7030 17377 7086
rect 17433 7030 17501 7086
rect 17557 7030 17625 7086
rect 17681 7030 17749 7086
rect 17805 7030 17907 7086
rect 17284 6962 17907 7030
rect 17284 6906 17377 6962
rect 17433 6906 17501 6962
rect 17557 6906 17625 6962
rect 17681 6906 17749 6962
rect 17805 6906 17907 6962
rect 17284 6838 17907 6906
rect 17284 6782 17377 6838
rect 17433 6782 17501 6838
rect 17557 6782 17625 6838
rect 17681 6782 17749 6838
rect 17805 6782 17907 6838
rect 17284 6714 17907 6782
rect 17284 6658 17377 6714
rect 17433 6658 17501 6714
rect 17557 6658 17625 6714
rect 17681 6658 17749 6714
rect 17805 6658 17907 6714
rect 17284 6590 17907 6658
rect 3953 6447 4017 6503
rect 4073 6447 4141 6503
rect 4197 6447 4265 6503
rect 4321 6447 4389 6503
rect 4445 6447 4513 6503
rect 4569 6447 4637 6503
rect 4693 6447 4761 6503
rect 4817 6447 4885 6503
rect 4941 6447 5009 6503
rect 5065 6447 5133 6503
rect 5189 6447 5257 6503
rect 5313 6447 5381 6503
rect 5437 6447 5505 6503
rect 5561 6447 5629 6503
rect 5685 6447 5753 6503
rect 5809 6447 5877 6503
rect 5933 6447 6001 6503
rect 6057 6447 6125 6503
rect 6181 6447 6249 6503
rect 6305 6447 6373 6503
rect 6429 6447 6493 6503
rect 3953 6379 6493 6447
rect 3953 6323 4017 6379
rect 4073 6323 4141 6379
rect 4197 6323 4265 6379
rect 4321 6323 4389 6379
rect 4445 6323 4513 6379
rect 4569 6323 4637 6379
rect 4693 6323 4761 6379
rect 4817 6323 4885 6379
rect 4941 6323 5009 6379
rect 5065 6323 5133 6379
rect 5189 6323 5257 6379
rect 5313 6323 5381 6379
rect 5437 6323 5505 6379
rect 5561 6323 5629 6379
rect 5685 6323 5753 6379
rect 5809 6323 5877 6379
rect 5933 6323 6001 6379
rect 6057 6323 6125 6379
rect 6181 6323 6249 6379
rect 6305 6323 6373 6379
rect 6429 6323 6493 6379
rect 3953 6255 6493 6323
rect 17284 6534 17377 6590
rect 17433 6534 17501 6590
rect 17557 6534 17625 6590
rect 17681 6534 17749 6590
rect 17805 6534 17907 6590
rect 17284 6466 17907 6534
rect 17284 6410 17377 6466
rect 17433 6410 17501 6466
rect 17557 6410 17625 6466
rect 17681 6410 17749 6466
rect 17805 6410 17907 6466
rect 17284 6306 17907 6410
rect 3953 6199 4017 6255
rect 4073 6199 4141 6255
rect 4197 6199 4265 6255
rect 4321 6199 4389 6255
rect 4445 6199 4513 6255
rect 4569 6199 4637 6255
rect 4693 6199 4761 6255
rect 4817 6199 4885 6255
rect 4941 6199 5009 6255
rect 5065 6199 5133 6255
rect 5189 6199 5257 6255
rect 5313 6199 5381 6255
rect 5437 6199 5505 6255
rect 5561 6199 5629 6255
rect 5685 6199 5753 6255
rect 5809 6199 5877 6255
rect 5933 6199 6001 6255
rect 6057 6199 6125 6255
rect 6181 6199 6249 6255
rect 6305 6199 6373 6255
rect 6429 6199 6493 6255
rect 3953 6131 6493 6199
rect 3953 6075 4017 6131
rect 4073 6075 4141 6131
rect 4197 6075 4265 6131
rect 4321 6075 4389 6131
rect 4445 6075 4513 6131
rect 4569 6075 4637 6131
rect 4693 6075 4761 6131
rect 4817 6075 4885 6131
rect 4941 6075 5009 6131
rect 5065 6075 5133 6131
rect 5189 6075 5257 6131
rect 5313 6075 5381 6131
rect 5437 6075 5505 6131
rect 5561 6075 5629 6131
rect 5685 6075 5753 6131
rect 5809 6075 5877 6131
rect 5933 6075 6001 6131
rect 6057 6075 6125 6131
rect 6181 6075 6249 6131
rect 6305 6075 6373 6131
rect 6429 6075 6493 6131
rect 3953 6007 6493 6075
rect 3953 5951 4017 6007
rect 4073 5951 4141 6007
rect 4197 5951 4265 6007
rect 4321 5951 4389 6007
rect 4445 5951 4513 6007
rect 4569 5951 4637 6007
rect 4693 5951 4761 6007
rect 4817 5951 4885 6007
rect 4941 5951 5009 6007
rect 5065 5951 5133 6007
rect 5189 5951 5257 6007
rect 5313 5951 5381 6007
rect 5437 5951 5505 6007
rect 5561 5951 5629 6007
rect 5685 5951 5753 6007
rect 5809 5951 5877 6007
rect 5933 5951 6001 6007
rect 6057 5951 6125 6007
rect 6181 5951 6249 6007
rect 6305 5951 6373 6007
rect 6429 5951 6493 6007
rect 3953 5884 6493 5951
<< via3 >>
rect 3977 8591 4033 8647
rect 4101 8591 4157 8647
rect 4225 8591 4281 8647
rect 4349 8591 4405 8647
rect 4473 8591 4529 8647
rect 4597 8591 4653 8647
rect 4721 8591 4777 8647
rect 4845 8591 4901 8647
rect 4969 8591 5025 8647
rect 5093 8591 5149 8647
rect 5217 8591 5273 8647
rect 5341 8591 5397 8647
rect 5465 8591 5521 8647
rect 5589 8591 5645 8647
rect 5713 8591 5769 8647
rect 5837 8591 5893 8647
rect 5961 8591 6017 8647
rect 6085 8591 6141 8647
rect 6209 8591 6265 8647
rect 6333 8591 6389 8647
rect 3977 8467 4033 8523
rect 4101 8467 4157 8523
rect 4225 8467 4281 8523
rect 4349 8467 4405 8523
rect 4473 8467 4529 8523
rect 4597 8467 4653 8523
rect 4721 8467 4777 8523
rect 4845 8467 4901 8523
rect 4969 8467 5025 8523
rect 5093 8467 5149 8523
rect 5217 8467 5273 8523
rect 5341 8467 5397 8523
rect 5465 8467 5521 8523
rect 5589 8467 5645 8523
rect 5713 8467 5769 8523
rect 5837 8467 5893 8523
rect 5961 8467 6017 8523
rect 6085 8467 6141 8523
rect 6209 8467 6265 8523
rect 6333 8467 6389 8523
rect 3977 8343 4033 8399
rect 4101 8343 4157 8399
rect 4225 8343 4281 8399
rect 4349 8343 4405 8399
rect 4473 8343 4529 8399
rect 4597 8343 4653 8399
rect 4721 8343 4777 8399
rect 4845 8343 4901 8399
rect 4969 8343 5025 8399
rect 5093 8343 5149 8399
rect 5217 8343 5273 8399
rect 5341 8343 5397 8399
rect 5465 8343 5521 8399
rect 5589 8343 5645 8399
rect 5713 8343 5769 8399
rect 5837 8343 5893 8399
rect 5961 8343 6017 8399
rect 6085 8343 6141 8399
rect 6209 8343 6265 8399
rect 6333 8343 6389 8399
rect 3977 8219 4033 8275
rect 4101 8219 4157 8275
rect 4225 8219 4281 8275
rect 4349 8219 4405 8275
rect 4473 8219 4529 8275
rect 4597 8219 4653 8275
rect 4721 8219 4777 8275
rect 4845 8219 4901 8275
rect 4969 8219 5025 8275
rect 5093 8219 5149 8275
rect 5217 8219 5273 8275
rect 5341 8219 5397 8275
rect 5465 8219 5521 8275
rect 5589 8219 5645 8275
rect 5713 8219 5769 8275
rect 5837 8219 5893 8275
rect 5961 8219 6017 8275
rect 6085 8219 6141 8275
rect 6209 8219 6265 8275
rect 6333 8219 6389 8275
rect 3977 8095 4033 8151
rect 4101 8095 4157 8151
rect 4225 8095 4281 8151
rect 4349 8095 4405 8151
rect 4473 8095 4529 8151
rect 4597 8095 4653 8151
rect 4721 8095 4777 8151
rect 4845 8095 4901 8151
rect 4969 8095 5025 8151
rect 5093 8095 5149 8151
rect 5217 8095 5273 8151
rect 5341 8095 5397 8151
rect 5465 8095 5521 8151
rect 5589 8095 5645 8151
rect 5713 8095 5769 8151
rect 5837 8095 5893 8151
rect 5961 8095 6017 8151
rect 6085 8095 6141 8151
rect 6209 8095 6265 8151
rect 6333 8095 6389 8151
rect 3977 7971 4033 8027
rect 4101 7971 4157 8027
rect 4225 7971 4281 8027
rect 4349 7971 4405 8027
rect 4473 7971 4529 8027
rect 4597 7971 4653 8027
rect 4721 7971 4777 8027
rect 4845 7971 4901 8027
rect 4969 7971 5025 8027
rect 5093 7971 5149 8027
rect 5217 7971 5273 8027
rect 5341 7971 5397 8027
rect 5465 7971 5521 8027
rect 5589 7971 5645 8027
rect 5713 7971 5769 8027
rect 5837 7971 5893 8027
rect 5961 7971 6017 8027
rect 6085 7971 6141 8027
rect 6209 7971 6265 8027
rect 6333 7971 6389 8027
rect 4017 6571 4073 6627
rect 4141 6571 4197 6627
rect 4265 6571 4321 6627
rect 4389 6571 4445 6627
rect 4513 6571 4569 6627
rect 4637 6571 4693 6627
rect 4761 6571 4817 6627
rect 4885 6571 4941 6627
rect 5009 6571 5065 6627
rect 5133 6571 5189 6627
rect 5257 6571 5313 6627
rect 5381 6571 5437 6627
rect 5505 6571 5561 6627
rect 5629 6571 5685 6627
rect 5753 6571 5809 6627
rect 5877 6571 5933 6627
rect 6001 6571 6057 6627
rect 6125 6571 6181 6627
rect 6249 6571 6305 6627
rect 6373 6571 6429 6627
rect 7093 6610 7199 7602
rect 7199 6610 7357 7602
rect 17377 7402 17433 7458
rect 17501 7402 17557 7458
rect 17625 7402 17681 7458
rect 17749 7402 17805 7458
rect 17377 7278 17433 7334
rect 17501 7278 17557 7334
rect 17625 7278 17681 7334
rect 17749 7278 17805 7334
rect 17377 7154 17433 7210
rect 17501 7154 17557 7210
rect 17625 7154 17681 7210
rect 17749 7154 17805 7210
rect 17377 7030 17433 7086
rect 17501 7030 17557 7086
rect 17625 7030 17681 7086
rect 17749 7030 17805 7086
rect 17377 6906 17433 6962
rect 17501 6906 17557 6962
rect 17625 6906 17681 6962
rect 17749 6906 17805 6962
rect 17377 6782 17433 6838
rect 17501 6782 17557 6838
rect 17625 6782 17681 6838
rect 17749 6782 17805 6838
rect 17377 6658 17433 6714
rect 17501 6658 17557 6714
rect 17625 6658 17681 6714
rect 17749 6658 17805 6714
rect 4017 6447 4073 6503
rect 4141 6447 4197 6503
rect 4265 6447 4321 6503
rect 4389 6447 4445 6503
rect 4513 6447 4569 6503
rect 4637 6447 4693 6503
rect 4761 6447 4817 6503
rect 4885 6447 4941 6503
rect 5009 6447 5065 6503
rect 5133 6447 5189 6503
rect 5257 6447 5313 6503
rect 5381 6447 5437 6503
rect 5505 6447 5561 6503
rect 5629 6447 5685 6503
rect 5753 6447 5809 6503
rect 5877 6447 5933 6503
rect 6001 6447 6057 6503
rect 6125 6447 6181 6503
rect 6249 6447 6305 6503
rect 6373 6447 6429 6503
rect 4017 6323 4073 6379
rect 4141 6323 4197 6379
rect 4265 6323 4321 6379
rect 4389 6323 4445 6379
rect 4513 6323 4569 6379
rect 4637 6323 4693 6379
rect 4761 6323 4817 6379
rect 4885 6323 4941 6379
rect 5009 6323 5065 6379
rect 5133 6323 5189 6379
rect 5257 6323 5313 6379
rect 5381 6323 5437 6379
rect 5505 6323 5561 6379
rect 5629 6323 5685 6379
rect 5753 6323 5809 6379
rect 5877 6323 5933 6379
rect 6001 6323 6057 6379
rect 6125 6323 6181 6379
rect 6249 6323 6305 6379
rect 6373 6323 6429 6379
rect 17377 6534 17433 6590
rect 17501 6534 17557 6590
rect 17625 6534 17681 6590
rect 17749 6534 17805 6590
rect 17377 6410 17433 6466
rect 17501 6410 17557 6466
rect 17625 6410 17681 6466
rect 17749 6410 17805 6466
rect 4017 6199 4073 6255
rect 4141 6199 4197 6255
rect 4265 6199 4321 6255
rect 4389 6199 4445 6255
rect 4513 6199 4569 6255
rect 4637 6199 4693 6255
rect 4761 6199 4817 6255
rect 4885 6199 4941 6255
rect 5009 6199 5065 6255
rect 5133 6199 5189 6255
rect 5257 6199 5313 6255
rect 5381 6199 5437 6255
rect 5505 6199 5561 6255
rect 5629 6199 5685 6255
rect 5753 6199 5809 6255
rect 5877 6199 5933 6255
rect 6001 6199 6057 6255
rect 6125 6199 6181 6255
rect 6249 6199 6305 6255
rect 6373 6199 6429 6255
rect 4017 6075 4073 6131
rect 4141 6075 4197 6131
rect 4265 6075 4321 6131
rect 4389 6075 4445 6131
rect 4513 6075 4569 6131
rect 4637 6075 4693 6131
rect 4761 6075 4817 6131
rect 4885 6075 4941 6131
rect 5009 6075 5065 6131
rect 5133 6075 5189 6131
rect 5257 6075 5313 6131
rect 5381 6075 5437 6131
rect 5505 6075 5561 6131
rect 5629 6075 5685 6131
rect 5753 6075 5809 6131
rect 5877 6075 5933 6131
rect 6001 6075 6057 6131
rect 6125 6075 6181 6131
rect 6249 6075 6305 6131
rect 6373 6075 6429 6131
rect 4017 5951 4073 6007
rect 4141 5951 4197 6007
rect 4265 5951 4321 6007
rect 4389 5951 4445 6007
rect 4513 5951 4569 6007
rect 4637 5951 4693 6007
rect 4761 5951 4817 6007
rect 4885 5951 4941 6007
rect 5009 5951 5065 6007
rect 5133 5951 5189 6007
rect 5257 5951 5313 6007
rect 5381 5951 5437 6007
rect 5505 5951 5561 6007
rect 5629 5951 5685 6007
rect 5753 5951 5809 6007
rect 5877 5951 5933 6007
rect 6001 5951 6057 6007
rect 6125 5951 6181 6007
rect 6249 5951 6305 6007
rect 6373 5951 6429 6007
<< metal4 >>
rect 3923 8647 6463 8714
rect 3923 8591 3977 8647
rect 4033 8591 4101 8647
rect 4157 8591 4225 8647
rect 4281 8591 4349 8647
rect 4405 8591 4473 8647
rect 4529 8591 4597 8647
rect 4653 8591 4721 8647
rect 4777 8591 4845 8647
rect 4901 8591 4969 8647
rect 5025 8591 5093 8647
rect 5149 8591 5217 8647
rect 5273 8591 5341 8647
rect 5397 8591 5465 8647
rect 5521 8591 5589 8647
rect 5645 8591 5713 8647
rect 5769 8591 5837 8647
rect 5893 8591 5961 8647
rect 6017 8591 6085 8647
rect 6141 8591 6209 8647
rect 6265 8591 6333 8647
rect 6389 8591 6463 8647
rect 3923 8523 6463 8591
rect 3923 8467 3977 8523
rect 4033 8467 4101 8523
rect 4157 8467 4225 8523
rect 4281 8467 4349 8523
rect 4405 8467 4473 8523
rect 4529 8467 4597 8523
rect 4653 8467 4721 8523
rect 4777 8467 4845 8523
rect 4901 8467 4969 8523
rect 5025 8467 5093 8523
rect 5149 8467 5217 8523
rect 5273 8467 5341 8523
rect 5397 8467 5465 8523
rect 5521 8467 5589 8523
rect 5645 8467 5713 8523
rect 5769 8467 5837 8523
rect 5893 8467 5961 8523
rect 6017 8467 6085 8523
rect 6141 8467 6209 8523
rect 6265 8467 6333 8523
rect 6389 8467 6463 8523
rect 3923 8399 6463 8467
rect 3923 8343 3977 8399
rect 4033 8343 4101 8399
rect 4157 8343 4225 8399
rect 4281 8343 4349 8399
rect 4405 8343 4473 8399
rect 4529 8343 4597 8399
rect 4653 8343 4721 8399
rect 4777 8343 4845 8399
rect 4901 8343 4969 8399
rect 5025 8343 5093 8399
rect 5149 8343 5217 8399
rect 5273 8343 5341 8399
rect 5397 8343 5465 8399
rect 5521 8343 5589 8399
rect 5645 8343 5713 8399
rect 5769 8343 5837 8399
rect 5893 8343 5961 8399
rect 6017 8343 6085 8399
rect 6141 8343 6209 8399
rect 6265 8343 6333 8399
rect 6389 8343 6463 8399
rect 3923 8275 6463 8343
rect 3923 8219 3977 8275
rect 4033 8219 4101 8275
rect 4157 8219 4225 8275
rect 4281 8219 4349 8275
rect 4405 8219 4473 8275
rect 4529 8219 4597 8275
rect 4653 8219 4721 8275
rect 4777 8219 4845 8275
rect 4901 8219 4969 8275
rect 5025 8219 5093 8275
rect 5149 8219 5217 8275
rect 5273 8219 5341 8275
rect 5397 8219 5465 8275
rect 5521 8219 5589 8275
rect 5645 8219 5713 8275
rect 5769 8219 5837 8275
rect 5893 8219 5961 8275
rect 6017 8219 6085 8275
rect 6141 8219 6209 8275
rect 6265 8219 6333 8275
rect 6389 8219 6463 8275
rect 3923 8151 6463 8219
rect 3923 8095 3977 8151
rect 4033 8095 4101 8151
rect 4157 8095 4225 8151
rect 4281 8095 4349 8151
rect 4405 8095 4473 8151
rect 4529 8095 4597 8151
rect 4653 8095 4721 8151
rect 4777 8095 4845 8151
rect 4901 8095 4969 8151
rect 5025 8095 5093 8151
rect 5149 8095 5217 8151
rect 5273 8095 5341 8151
rect 5397 8095 5465 8151
rect 5521 8095 5589 8151
rect 5645 8095 5713 8151
rect 5769 8095 5837 8151
rect 5893 8095 5961 8151
rect 6017 8095 6085 8151
rect 6141 8095 6209 8151
rect 6265 8095 6333 8151
rect 6389 8095 6463 8151
rect 3923 8027 6463 8095
rect 3923 7971 3977 8027
rect 4033 7971 4101 8027
rect 4157 7971 4225 8027
rect 4281 7971 4349 8027
rect 4405 7971 4473 8027
rect 4529 7971 4597 8027
rect 4653 7971 4721 8027
rect 4777 7971 4845 8027
rect 4901 7971 4969 8027
rect 5025 7971 5093 8027
rect 5149 7971 5217 8027
rect 5273 7971 5341 8027
rect 5397 7971 5465 8027
rect 5521 7971 5589 8027
rect 5645 7971 5713 8027
rect 5769 7971 5837 8027
rect 5893 7971 5961 8027
rect 6017 7971 6085 8027
rect 6141 7971 6209 8027
rect 6265 7971 6333 8027
rect 6389 7971 6463 8027
rect 3923 7914 6463 7971
rect 7046 7602 7414 7647
rect 3953 6627 6493 6684
rect 3953 6571 4017 6627
rect 4073 6571 4141 6627
rect 4197 6571 4265 6627
rect 4321 6571 4389 6627
rect 4445 6571 4513 6627
rect 4569 6571 4637 6627
rect 4693 6571 4761 6627
rect 4817 6571 4885 6627
rect 4941 6571 5009 6627
rect 5065 6571 5133 6627
rect 5189 6571 5257 6627
rect 5313 6571 5381 6627
rect 5437 6571 5505 6627
rect 5561 6571 5629 6627
rect 5685 6571 5753 6627
rect 5809 6571 5877 6627
rect 5933 6571 6001 6627
rect 6057 6571 6125 6627
rect 6181 6571 6249 6627
rect 6305 6571 6373 6627
rect 6429 6571 6493 6627
rect 3953 6503 6493 6571
rect 7046 6610 7093 7602
rect 7357 6610 7414 7602
rect 17284 7458 17907 7555
rect 17284 7402 17377 7458
rect 17433 7402 17501 7458
rect 17557 7402 17625 7458
rect 17681 7402 17749 7458
rect 17805 7402 17907 7458
rect 17284 7334 17907 7402
rect 17284 7278 17377 7334
rect 17433 7278 17501 7334
rect 17557 7278 17625 7334
rect 17681 7278 17749 7334
rect 17805 7278 17907 7334
rect 7046 6561 7414 6610
rect 15694 7184 17016 7256
rect 15694 7128 15826 7184
rect 15882 7128 15950 7184
rect 16006 7128 16074 7184
rect 16130 7128 16198 7184
rect 16254 7128 16322 7184
rect 16378 7128 16446 7184
rect 16502 7128 16570 7184
rect 16626 7128 16694 7184
rect 16750 7128 16818 7184
rect 16874 7128 17016 7184
rect 15694 7060 17016 7128
rect 15694 7004 15826 7060
rect 15882 7004 15950 7060
rect 16006 7004 16074 7060
rect 16130 7004 16198 7060
rect 16254 7004 16322 7060
rect 16378 7004 16446 7060
rect 16502 7004 16570 7060
rect 16626 7004 16694 7060
rect 16750 7004 16818 7060
rect 16874 7004 17016 7060
rect 15694 6936 17016 7004
rect 15694 6880 15826 6936
rect 15882 6880 15950 6936
rect 16006 6880 16074 6936
rect 16130 6880 16198 6936
rect 16254 6880 16322 6936
rect 16378 6880 16446 6936
rect 16502 6880 16570 6936
rect 16626 6880 16694 6936
rect 16750 6880 16818 6936
rect 16874 6880 17016 6936
rect 15694 6812 17016 6880
rect 15694 6756 15826 6812
rect 15882 6756 15950 6812
rect 16006 6756 16074 6812
rect 16130 6756 16198 6812
rect 16254 6756 16322 6812
rect 16378 6756 16446 6812
rect 16502 6756 16570 6812
rect 16626 6756 16694 6812
rect 16750 6756 16818 6812
rect 16874 6756 17016 6812
rect 15694 6688 17016 6756
rect 15694 6632 15826 6688
rect 15882 6632 15950 6688
rect 16006 6632 16074 6688
rect 16130 6632 16198 6688
rect 16254 6632 16322 6688
rect 16378 6632 16446 6688
rect 16502 6632 16570 6688
rect 16626 6632 16694 6688
rect 16750 6632 16818 6688
rect 16874 6632 17016 6688
rect 15694 6564 17016 6632
rect 3953 6447 4017 6503
rect 4073 6447 4141 6503
rect 4197 6447 4265 6503
rect 4321 6447 4389 6503
rect 4445 6447 4513 6503
rect 4569 6447 4637 6503
rect 4693 6447 4761 6503
rect 4817 6447 4885 6503
rect 4941 6447 5009 6503
rect 5065 6447 5133 6503
rect 5189 6447 5257 6503
rect 5313 6447 5381 6503
rect 5437 6447 5505 6503
rect 5561 6447 5629 6503
rect 5685 6447 5753 6503
rect 5809 6447 5877 6503
rect 5933 6447 6001 6503
rect 6057 6447 6125 6503
rect 6181 6447 6249 6503
rect 6305 6447 6373 6503
rect 6429 6447 6493 6503
rect 3953 6379 6493 6447
rect 3953 6323 4017 6379
rect 4073 6323 4141 6379
rect 4197 6323 4265 6379
rect 4321 6323 4389 6379
rect 4445 6323 4513 6379
rect 4569 6323 4637 6379
rect 4693 6323 4761 6379
rect 4817 6323 4885 6379
rect 4941 6323 5009 6379
rect 5065 6323 5133 6379
rect 5189 6323 5257 6379
rect 5313 6323 5381 6379
rect 5437 6323 5505 6379
rect 5561 6323 5629 6379
rect 5685 6323 5753 6379
rect 5809 6323 5877 6379
rect 5933 6323 6001 6379
rect 6057 6323 6125 6379
rect 6181 6323 6249 6379
rect 6305 6323 6373 6379
rect 6429 6323 6493 6379
rect 3953 6255 6493 6323
rect 3953 6199 4017 6255
rect 4073 6199 4141 6255
rect 4197 6199 4265 6255
rect 4321 6199 4389 6255
rect 4445 6199 4513 6255
rect 4569 6199 4637 6255
rect 4693 6199 4761 6255
rect 4817 6199 4885 6255
rect 4941 6199 5009 6255
rect 5065 6199 5133 6255
rect 5189 6199 5257 6255
rect 5313 6199 5381 6255
rect 5437 6199 5505 6255
rect 5561 6199 5629 6255
rect 5685 6199 5753 6255
rect 5809 6199 5877 6255
rect 5933 6199 6001 6255
rect 6057 6199 6125 6255
rect 6181 6199 6249 6255
rect 6305 6199 6373 6255
rect 6429 6199 6493 6255
rect 3953 6131 6493 6199
rect 3953 6075 4017 6131
rect 4073 6075 4141 6131
rect 4197 6075 4265 6131
rect 4321 6075 4389 6131
rect 4445 6075 4513 6131
rect 4569 6075 4637 6131
rect 4693 6075 4761 6131
rect 4817 6075 4885 6131
rect 4941 6075 5009 6131
rect 5065 6075 5133 6131
rect 5189 6075 5257 6131
rect 5313 6075 5381 6131
rect 5437 6075 5505 6131
rect 5561 6075 5629 6131
rect 5685 6075 5753 6131
rect 5809 6075 5877 6131
rect 5933 6075 6001 6131
rect 6057 6075 6125 6131
rect 6181 6075 6249 6131
rect 6305 6075 6373 6131
rect 6429 6075 6493 6131
rect 3953 6007 6493 6075
rect 3953 5951 4017 6007
rect 4073 5951 4141 6007
rect 4197 5951 4265 6007
rect 4321 5951 4389 6007
rect 4445 5951 4513 6007
rect 4569 5951 4637 6007
rect 4693 5951 4761 6007
rect 4817 5951 4885 6007
rect 4941 5951 5009 6007
rect 5065 5951 5133 6007
rect 5189 5951 5257 6007
rect 5313 5951 5381 6007
rect 5437 5951 5505 6007
rect 5561 5951 5629 6007
rect 5685 5951 5753 6007
rect 5809 5951 5877 6007
rect 5933 5951 6001 6007
rect 6057 5951 6125 6007
rect 6181 5951 6249 6007
rect 6305 5951 6373 6007
rect 6429 5951 6493 6007
rect 3953 5884 6493 5951
rect 15694 6508 15826 6564
rect 15882 6508 15950 6564
rect 16006 6508 16074 6564
rect 16130 6508 16198 6564
rect 16254 6508 16322 6564
rect 16378 6508 16446 6564
rect 16502 6508 16570 6564
rect 16626 6508 16694 6564
rect 16750 6508 16818 6564
rect 16874 6508 17016 6564
rect 15694 6440 17016 6508
rect 15694 6384 15826 6440
rect 15882 6384 15950 6440
rect 16006 6384 16074 6440
rect 16130 6384 16198 6440
rect 16254 6384 16322 6440
rect 16378 6384 16446 6440
rect 16502 6384 16570 6440
rect 16626 6384 16694 6440
rect 16750 6384 16818 6440
rect 16874 6384 17016 6440
rect 15694 6316 17016 6384
rect 15694 6260 15826 6316
rect 15882 6260 15950 6316
rect 16006 6260 16074 6316
rect 16130 6260 16198 6316
rect 16254 6260 16322 6316
rect 16378 6260 16446 6316
rect 16502 6260 16570 6316
rect 16626 6260 16694 6316
rect 16750 6260 16818 6316
rect 16874 6260 17016 6316
rect 17284 7210 17907 7278
rect 17284 7154 17377 7210
rect 17433 7154 17501 7210
rect 17557 7154 17625 7210
rect 17681 7154 17749 7210
rect 17805 7154 17907 7210
rect 17284 7086 17907 7154
rect 17284 7030 17377 7086
rect 17433 7030 17501 7086
rect 17557 7030 17625 7086
rect 17681 7030 17749 7086
rect 17805 7030 17907 7086
rect 17284 6962 17907 7030
rect 17284 6906 17377 6962
rect 17433 6906 17501 6962
rect 17557 6906 17625 6962
rect 17681 6906 17749 6962
rect 17805 6906 17907 6962
rect 17284 6838 17907 6906
rect 17284 6782 17377 6838
rect 17433 6782 17501 6838
rect 17557 6782 17625 6838
rect 17681 6782 17749 6838
rect 17805 6782 17907 6838
rect 17284 6714 17907 6782
rect 17284 6658 17377 6714
rect 17433 6658 17501 6714
rect 17557 6658 17625 6714
rect 17681 6658 17749 6714
rect 17805 6658 17907 6714
rect 17284 6590 17907 6658
rect 17284 6534 17377 6590
rect 17433 6534 17501 6590
rect 17557 6534 17625 6590
rect 17681 6534 17749 6590
rect 17805 6534 17907 6590
rect 17284 6466 17907 6534
rect 17284 6410 17377 6466
rect 17433 6410 17501 6466
rect 17557 6410 17625 6466
rect 17681 6410 17749 6466
rect 17805 6410 17907 6466
rect 17284 6306 17907 6410
rect 15694 6192 17016 6260
rect 15694 6136 15826 6192
rect 15882 6136 15950 6192
rect 16006 6136 16074 6192
rect 16130 6136 16198 6192
rect 16254 6136 16322 6192
rect 16378 6136 16446 6192
rect 16502 6136 16570 6192
rect 16626 6136 16694 6192
rect 16750 6136 16818 6192
rect 16874 6136 17016 6192
rect 15694 6068 17016 6136
rect 15694 6012 15826 6068
rect 15882 6012 15950 6068
rect 16006 6012 16074 6068
rect 16130 6012 16198 6068
rect 16254 6012 16322 6068
rect 16378 6012 16446 6068
rect 16502 6012 16570 6068
rect 16626 6012 16694 6068
rect 16750 6012 16818 6068
rect 16874 6012 17016 6068
rect 15694 5944 17016 6012
rect 15694 5888 15826 5944
rect 15882 5888 15950 5944
rect 16006 5888 16074 5944
rect 16130 5888 16198 5944
rect 16254 5888 16322 5944
rect 16378 5888 16446 5944
rect 16502 5888 16570 5944
rect 16626 5888 16694 5944
rect 16750 5888 16818 5944
rect 16874 5888 17016 5944
rect 15694 5808 17016 5888
<< via4 >>
rect 3977 8591 4033 8647
rect 4101 8591 4157 8647
rect 4225 8591 4281 8647
rect 4349 8591 4405 8647
rect 4473 8591 4529 8647
rect 4597 8591 4653 8647
rect 4721 8591 4777 8647
rect 4845 8591 4901 8647
rect 4969 8591 5025 8647
rect 5093 8591 5149 8647
rect 5217 8591 5273 8647
rect 5341 8591 5397 8647
rect 5465 8591 5521 8647
rect 5589 8591 5645 8647
rect 5713 8591 5769 8647
rect 5837 8591 5893 8647
rect 5961 8591 6017 8647
rect 6085 8591 6141 8647
rect 6209 8591 6265 8647
rect 6333 8591 6389 8647
rect 3977 8467 4033 8523
rect 4101 8467 4157 8523
rect 4225 8467 4281 8523
rect 4349 8467 4405 8523
rect 4473 8467 4529 8523
rect 4597 8467 4653 8523
rect 4721 8467 4777 8523
rect 4845 8467 4901 8523
rect 4969 8467 5025 8523
rect 5093 8467 5149 8523
rect 5217 8467 5273 8523
rect 5341 8467 5397 8523
rect 5465 8467 5521 8523
rect 5589 8467 5645 8523
rect 5713 8467 5769 8523
rect 5837 8467 5893 8523
rect 5961 8467 6017 8523
rect 6085 8467 6141 8523
rect 6209 8467 6265 8523
rect 6333 8467 6389 8523
rect 3977 8343 4033 8399
rect 4101 8343 4157 8399
rect 4225 8343 4281 8399
rect 4349 8343 4405 8399
rect 4473 8343 4529 8399
rect 4597 8343 4653 8399
rect 4721 8343 4777 8399
rect 4845 8343 4901 8399
rect 4969 8343 5025 8399
rect 5093 8343 5149 8399
rect 5217 8343 5273 8399
rect 5341 8343 5397 8399
rect 5465 8343 5521 8399
rect 5589 8343 5645 8399
rect 5713 8343 5769 8399
rect 5837 8343 5893 8399
rect 5961 8343 6017 8399
rect 6085 8343 6141 8399
rect 6209 8343 6265 8399
rect 6333 8343 6389 8399
rect 3977 8219 4033 8275
rect 4101 8219 4157 8275
rect 4225 8219 4281 8275
rect 4349 8219 4405 8275
rect 4473 8219 4529 8275
rect 4597 8219 4653 8275
rect 4721 8219 4777 8275
rect 4845 8219 4901 8275
rect 4969 8219 5025 8275
rect 5093 8219 5149 8275
rect 5217 8219 5273 8275
rect 5341 8219 5397 8275
rect 5465 8219 5521 8275
rect 5589 8219 5645 8275
rect 5713 8219 5769 8275
rect 5837 8219 5893 8275
rect 5961 8219 6017 8275
rect 6085 8219 6141 8275
rect 6209 8219 6265 8275
rect 6333 8219 6389 8275
rect 3977 8095 4033 8151
rect 4101 8095 4157 8151
rect 4225 8095 4281 8151
rect 4349 8095 4405 8151
rect 4473 8095 4529 8151
rect 4597 8095 4653 8151
rect 4721 8095 4777 8151
rect 4845 8095 4901 8151
rect 4969 8095 5025 8151
rect 5093 8095 5149 8151
rect 5217 8095 5273 8151
rect 5341 8095 5397 8151
rect 5465 8095 5521 8151
rect 5589 8095 5645 8151
rect 5713 8095 5769 8151
rect 5837 8095 5893 8151
rect 5961 8095 6017 8151
rect 6085 8095 6141 8151
rect 6209 8095 6265 8151
rect 6333 8095 6389 8151
rect 3977 7971 4033 8027
rect 4101 7971 4157 8027
rect 4225 7971 4281 8027
rect 4349 7971 4405 8027
rect 4473 7971 4529 8027
rect 4597 7971 4653 8027
rect 4721 7971 4777 8027
rect 4845 7971 4901 8027
rect 4969 7971 5025 8027
rect 5093 7971 5149 8027
rect 5217 7971 5273 8027
rect 5341 7971 5397 8027
rect 5465 7971 5521 8027
rect 5589 7971 5645 8027
rect 5713 7971 5769 8027
rect 5837 7971 5893 8027
rect 5961 7971 6017 8027
rect 6085 7971 6141 8027
rect 6209 7971 6265 8027
rect 6333 7971 6389 8027
rect 4017 6571 4073 6627
rect 4141 6571 4197 6627
rect 4265 6571 4321 6627
rect 4389 6571 4445 6627
rect 4513 6571 4569 6627
rect 4637 6571 4693 6627
rect 4761 6571 4817 6627
rect 4885 6571 4941 6627
rect 5009 6571 5065 6627
rect 5133 6571 5189 6627
rect 5257 6571 5313 6627
rect 5381 6571 5437 6627
rect 5505 6571 5561 6627
rect 5629 6571 5685 6627
rect 5753 6571 5809 6627
rect 5877 6571 5933 6627
rect 6001 6571 6057 6627
rect 6125 6571 6181 6627
rect 6249 6571 6305 6627
rect 6373 6571 6429 6627
rect 7093 6610 7357 7602
rect 17377 7402 17433 7458
rect 17501 7402 17557 7458
rect 17625 7402 17681 7458
rect 17749 7402 17805 7458
rect 17377 7278 17433 7334
rect 17501 7278 17557 7334
rect 17625 7278 17681 7334
rect 17749 7278 17805 7334
rect 15826 7128 15882 7184
rect 15950 7128 16006 7184
rect 16074 7128 16130 7184
rect 16198 7128 16254 7184
rect 16322 7128 16378 7184
rect 16446 7128 16502 7184
rect 16570 7128 16626 7184
rect 16694 7128 16750 7184
rect 16818 7128 16874 7184
rect 15826 7004 15882 7060
rect 15950 7004 16006 7060
rect 16074 7004 16130 7060
rect 16198 7004 16254 7060
rect 16322 7004 16378 7060
rect 16446 7004 16502 7060
rect 16570 7004 16626 7060
rect 16694 7004 16750 7060
rect 16818 7004 16874 7060
rect 15826 6880 15882 6936
rect 15950 6880 16006 6936
rect 16074 6880 16130 6936
rect 16198 6880 16254 6936
rect 16322 6880 16378 6936
rect 16446 6880 16502 6936
rect 16570 6880 16626 6936
rect 16694 6880 16750 6936
rect 16818 6880 16874 6936
rect 15826 6756 15882 6812
rect 15950 6756 16006 6812
rect 16074 6756 16130 6812
rect 16198 6756 16254 6812
rect 16322 6756 16378 6812
rect 16446 6756 16502 6812
rect 16570 6756 16626 6812
rect 16694 6756 16750 6812
rect 16818 6756 16874 6812
rect 15826 6632 15882 6688
rect 15950 6632 16006 6688
rect 16074 6632 16130 6688
rect 16198 6632 16254 6688
rect 16322 6632 16378 6688
rect 16446 6632 16502 6688
rect 16570 6632 16626 6688
rect 16694 6632 16750 6688
rect 16818 6632 16874 6688
rect 4017 6447 4073 6503
rect 4141 6447 4197 6503
rect 4265 6447 4321 6503
rect 4389 6447 4445 6503
rect 4513 6447 4569 6503
rect 4637 6447 4693 6503
rect 4761 6447 4817 6503
rect 4885 6447 4941 6503
rect 5009 6447 5065 6503
rect 5133 6447 5189 6503
rect 5257 6447 5313 6503
rect 5381 6447 5437 6503
rect 5505 6447 5561 6503
rect 5629 6447 5685 6503
rect 5753 6447 5809 6503
rect 5877 6447 5933 6503
rect 6001 6447 6057 6503
rect 6125 6447 6181 6503
rect 6249 6447 6305 6503
rect 6373 6447 6429 6503
rect 4017 6323 4073 6379
rect 4141 6323 4197 6379
rect 4265 6323 4321 6379
rect 4389 6323 4445 6379
rect 4513 6323 4569 6379
rect 4637 6323 4693 6379
rect 4761 6323 4817 6379
rect 4885 6323 4941 6379
rect 5009 6323 5065 6379
rect 5133 6323 5189 6379
rect 5257 6323 5313 6379
rect 5381 6323 5437 6379
rect 5505 6323 5561 6379
rect 5629 6323 5685 6379
rect 5753 6323 5809 6379
rect 5877 6323 5933 6379
rect 6001 6323 6057 6379
rect 6125 6323 6181 6379
rect 6249 6323 6305 6379
rect 6373 6323 6429 6379
rect 4017 6199 4073 6255
rect 4141 6199 4197 6255
rect 4265 6199 4321 6255
rect 4389 6199 4445 6255
rect 4513 6199 4569 6255
rect 4637 6199 4693 6255
rect 4761 6199 4817 6255
rect 4885 6199 4941 6255
rect 5009 6199 5065 6255
rect 5133 6199 5189 6255
rect 5257 6199 5313 6255
rect 5381 6199 5437 6255
rect 5505 6199 5561 6255
rect 5629 6199 5685 6255
rect 5753 6199 5809 6255
rect 5877 6199 5933 6255
rect 6001 6199 6057 6255
rect 6125 6199 6181 6255
rect 6249 6199 6305 6255
rect 6373 6199 6429 6255
rect 4017 6075 4073 6131
rect 4141 6075 4197 6131
rect 4265 6075 4321 6131
rect 4389 6075 4445 6131
rect 4513 6075 4569 6131
rect 4637 6075 4693 6131
rect 4761 6075 4817 6131
rect 4885 6075 4941 6131
rect 5009 6075 5065 6131
rect 5133 6075 5189 6131
rect 5257 6075 5313 6131
rect 5381 6075 5437 6131
rect 5505 6075 5561 6131
rect 5629 6075 5685 6131
rect 5753 6075 5809 6131
rect 5877 6075 5933 6131
rect 6001 6075 6057 6131
rect 6125 6075 6181 6131
rect 6249 6075 6305 6131
rect 6373 6075 6429 6131
rect 4017 5951 4073 6007
rect 4141 5951 4197 6007
rect 4265 5951 4321 6007
rect 4389 5951 4445 6007
rect 4513 5951 4569 6007
rect 4637 5951 4693 6007
rect 4761 5951 4817 6007
rect 4885 5951 4941 6007
rect 5009 5951 5065 6007
rect 5133 5951 5189 6007
rect 5257 5951 5313 6007
rect 5381 5951 5437 6007
rect 5505 5951 5561 6007
rect 5629 5951 5685 6007
rect 5753 5951 5809 6007
rect 5877 5951 5933 6007
rect 6001 5951 6057 6007
rect 6125 5951 6181 6007
rect 6249 5951 6305 6007
rect 6373 5951 6429 6007
rect 15826 6508 15882 6564
rect 15950 6508 16006 6564
rect 16074 6508 16130 6564
rect 16198 6508 16254 6564
rect 16322 6508 16378 6564
rect 16446 6508 16502 6564
rect 16570 6508 16626 6564
rect 16694 6508 16750 6564
rect 16818 6508 16874 6564
rect 15826 6384 15882 6440
rect 15950 6384 16006 6440
rect 16074 6384 16130 6440
rect 16198 6384 16254 6440
rect 16322 6384 16378 6440
rect 16446 6384 16502 6440
rect 16570 6384 16626 6440
rect 16694 6384 16750 6440
rect 16818 6384 16874 6440
rect 15826 6260 15882 6316
rect 15950 6260 16006 6316
rect 16074 6260 16130 6316
rect 16198 6260 16254 6316
rect 16322 6260 16378 6316
rect 16446 6260 16502 6316
rect 16570 6260 16626 6316
rect 16694 6260 16750 6316
rect 16818 6260 16874 6316
rect 17377 7154 17433 7210
rect 17501 7154 17557 7210
rect 17625 7154 17681 7210
rect 17749 7154 17805 7210
rect 17377 7030 17433 7086
rect 17501 7030 17557 7086
rect 17625 7030 17681 7086
rect 17749 7030 17805 7086
rect 17377 6906 17433 6962
rect 17501 6906 17557 6962
rect 17625 6906 17681 6962
rect 17749 6906 17805 6962
rect 17377 6782 17433 6838
rect 17501 6782 17557 6838
rect 17625 6782 17681 6838
rect 17749 6782 17805 6838
rect 17377 6658 17433 6714
rect 17501 6658 17557 6714
rect 17625 6658 17681 6714
rect 17749 6658 17805 6714
rect 17377 6534 17433 6590
rect 17501 6534 17557 6590
rect 17625 6534 17681 6590
rect 17749 6534 17805 6590
rect 17377 6410 17433 6466
rect 17501 6410 17557 6466
rect 17625 6410 17681 6466
rect 17749 6410 17805 6466
rect 15826 6136 15882 6192
rect 15950 6136 16006 6192
rect 16074 6136 16130 6192
rect 16198 6136 16254 6192
rect 16322 6136 16378 6192
rect 16446 6136 16502 6192
rect 16570 6136 16626 6192
rect 16694 6136 16750 6192
rect 16818 6136 16874 6192
rect 15826 6012 15882 6068
rect 15950 6012 16006 6068
rect 16074 6012 16130 6068
rect 16198 6012 16254 6068
rect 16322 6012 16378 6068
rect 16446 6012 16502 6068
rect 16570 6012 16626 6068
rect 16694 6012 16750 6068
rect 16818 6012 16874 6068
rect 15826 5888 15882 5944
rect 15950 5888 16006 5944
rect 16074 5888 16130 5944
rect 16198 5888 16254 5944
rect 16322 5888 16378 5944
rect 16446 5888 16502 5944
rect 16570 5888 16626 5944
rect 16694 5888 16750 5944
rect 16818 5888 16874 5944
<< metal5 >>
rect 24 8647 6463 8714
rect 24 8591 3977 8647
rect 4033 8591 4101 8647
rect 4157 8591 4225 8647
rect 4281 8591 4349 8647
rect 4405 8591 4473 8647
rect 4529 8591 4597 8647
rect 4653 8591 4721 8647
rect 4777 8591 4845 8647
rect 4901 8591 4969 8647
rect 5025 8591 5093 8647
rect 5149 8591 5217 8647
rect 5273 8591 5341 8647
rect 5397 8591 5465 8647
rect 5521 8591 5589 8647
rect 5645 8591 5713 8647
rect 5769 8591 5837 8647
rect 5893 8591 5961 8647
rect 6017 8591 6085 8647
rect 6141 8591 6209 8647
rect 6265 8591 6333 8647
rect 6389 8591 6463 8647
rect 24 8523 6463 8591
rect 24 8467 3977 8523
rect 4033 8467 4101 8523
rect 4157 8467 4225 8523
rect 4281 8467 4349 8523
rect 4405 8467 4473 8523
rect 4529 8467 4597 8523
rect 4653 8467 4721 8523
rect 4777 8467 4845 8523
rect 4901 8467 4969 8523
rect 5025 8467 5093 8523
rect 5149 8467 5217 8523
rect 5273 8467 5341 8523
rect 5397 8467 5465 8523
rect 5521 8467 5589 8523
rect 5645 8467 5713 8523
rect 5769 8467 5837 8523
rect 5893 8467 5961 8523
rect 6017 8467 6085 8523
rect 6141 8467 6209 8523
rect 6265 8467 6333 8523
rect 6389 8467 6463 8523
rect 24 8399 6463 8467
rect 24 8343 3977 8399
rect 4033 8343 4101 8399
rect 4157 8343 4225 8399
rect 4281 8343 4349 8399
rect 4405 8343 4473 8399
rect 4529 8343 4597 8399
rect 4653 8343 4721 8399
rect 4777 8343 4845 8399
rect 4901 8343 4969 8399
rect 5025 8343 5093 8399
rect 5149 8343 5217 8399
rect 5273 8343 5341 8399
rect 5397 8343 5465 8399
rect 5521 8343 5589 8399
rect 5645 8343 5713 8399
rect 5769 8343 5837 8399
rect 5893 8343 5961 8399
rect 6017 8343 6085 8399
rect 6141 8343 6209 8399
rect 6265 8343 6333 8399
rect 6389 8343 6463 8399
rect 24 8275 6463 8343
rect 24 8219 3977 8275
rect 4033 8219 4101 8275
rect 4157 8219 4225 8275
rect 4281 8219 4349 8275
rect 4405 8219 4473 8275
rect 4529 8219 4597 8275
rect 4653 8219 4721 8275
rect 4777 8219 4845 8275
rect 4901 8219 4969 8275
rect 5025 8219 5093 8275
rect 5149 8219 5217 8275
rect 5273 8219 5341 8275
rect 5397 8219 5465 8275
rect 5521 8219 5589 8275
rect 5645 8219 5713 8275
rect 5769 8219 5837 8275
rect 5893 8219 5961 8275
rect 6017 8219 6085 8275
rect 6141 8219 6209 8275
rect 6265 8219 6333 8275
rect 6389 8219 6463 8275
rect 24 8151 6463 8219
rect 24 8095 3977 8151
rect 4033 8095 4101 8151
rect 4157 8095 4225 8151
rect 4281 8095 4349 8151
rect 4405 8095 4473 8151
rect 4529 8095 4597 8151
rect 4653 8095 4721 8151
rect 4777 8095 4845 8151
rect 4901 8095 4969 8151
rect 5025 8095 5093 8151
rect 5149 8095 5217 8151
rect 5273 8095 5341 8151
rect 5397 8095 5465 8151
rect 5521 8095 5589 8151
rect 5645 8095 5713 8151
rect 5769 8095 5837 8151
rect 5893 8095 5961 8151
rect 6017 8095 6085 8151
rect 6141 8095 6209 8151
rect 6265 8095 6333 8151
rect 6389 8095 6463 8151
rect 24 8027 6463 8095
rect 24 7971 3977 8027
rect 4033 7971 4101 8027
rect 4157 7971 4225 8027
rect 4281 7971 4349 8027
rect 4405 7971 4473 8027
rect 4529 7971 4597 8027
rect 4653 7971 4721 8027
rect 4777 7971 4845 8027
rect 4901 7971 4969 8027
rect 5025 7971 5093 8027
rect 5149 7971 5217 8027
rect 5273 7971 5341 8027
rect 5397 7971 5465 8027
rect 5521 7971 5589 8027
rect 5645 7971 5713 8027
rect 5769 7971 5837 8027
rect 5893 7971 5961 8027
rect 6017 7971 6085 8027
rect 6141 7971 6209 8027
rect 6265 7971 6333 8027
rect 6389 7971 6463 8027
rect 24 7914 6463 7971
rect 7157 7735 17700 7983
rect 7157 7647 7414 7735
rect 7046 7602 7414 7647
rect 24 6627 6493 6684
rect 24 6571 4017 6627
rect 4073 6571 4141 6627
rect 4197 6571 4265 6627
rect 4321 6571 4389 6627
rect 4445 6571 4513 6627
rect 4569 6571 4637 6627
rect 4693 6571 4761 6627
rect 4817 6571 4885 6627
rect 4941 6571 5009 6627
rect 5065 6571 5133 6627
rect 5189 6571 5257 6627
rect 5313 6571 5381 6627
rect 5437 6571 5505 6627
rect 5561 6571 5629 6627
rect 5685 6571 5753 6627
rect 5809 6571 5877 6627
rect 5933 6571 6001 6627
rect 6057 6571 6125 6627
rect 6181 6571 6249 6627
rect 6305 6571 6373 6627
rect 6429 6571 6493 6627
rect 24 6503 6493 6571
rect 7046 6610 7093 7602
rect 7357 6610 7414 7602
rect 17284 7619 17700 7735
rect 17284 7458 17907 7619
rect 17284 7402 17377 7458
rect 17433 7402 17501 7458
rect 17557 7402 17625 7458
rect 17681 7402 17749 7458
rect 17805 7402 17907 7458
rect 17284 7334 17907 7402
rect 17284 7278 17377 7334
rect 17433 7278 17501 7334
rect 17557 7278 17625 7334
rect 17681 7278 17749 7334
rect 17805 7278 17907 7334
rect 7046 6561 7414 6610
rect 15454 7184 17016 7256
rect 15454 7128 15826 7184
rect 15882 7128 15950 7184
rect 16006 7128 16074 7184
rect 16130 7128 16198 7184
rect 16254 7128 16322 7184
rect 16378 7128 16446 7184
rect 16502 7128 16570 7184
rect 16626 7128 16694 7184
rect 16750 7128 16818 7184
rect 16874 7128 17016 7184
rect 15454 7060 17016 7128
rect 15454 7004 15826 7060
rect 15882 7004 15950 7060
rect 16006 7004 16074 7060
rect 16130 7004 16198 7060
rect 16254 7004 16322 7060
rect 16378 7004 16446 7060
rect 16502 7004 16570 7060
rect 16626 7004 16694 7060
rect 16750 7004 16818 7060
rect 16874 7004 17016 7060
rect 15454 6936 17016 7004
rect 15454 6880 15826 6936
rect 15882 6880 15950 6936
rect 16006 6880 16074 6936
rect 16130 6880 16198 6936
rect 16254 6880 16322 6936
rect 16378 6880 16446 6936
rect 16502 6880 16570 6936
rect 16626 6880 16694 6936
rect 16750 6880 16818 6936
rect 16874 6880 17016 6936
rect 15454 6812 17016 6880
rect 15454 6756 15826 6812
rect 15882 6756 15950 6812
rect 16006 6756 16074 6812
rect 16130 6756 16198 6812
rect 16254 6756 16322 6812
rect 16378 6756 16446 6812
rect 16502 6756 16570 6812
rect 16626 6756 16694 6812
rect 16750 6756 16818 6812
rect 16874 6756 17016 6812
rect 15454 6688 17016 6756
rect 15454 6632 15826 6688
rect 15882 6632 15950 6688
rect 16006 6632 16074 6688
rect 16130 6632 16198 6688
rect 16254 6632 16322 6688
rect 16378 6632 16446 6688
rect 16502 6632 16570 6688
rect 16626 6632 16694 6688
rect 16750 6632 16818 6688
rect 16874 6632 17016 6688
rect 15454 6564 17016 6632
rect 24 6447 4017 6503
rect 4073 6447 4141 6503
rect 4197 6447 4265 6503
rect 4321 6447 4389 6503
rect 4445 6447 4513 6503
rect 4569 6447 4637 6503
rect 4693 6447 4761 6503
rect 4817 6447 4885 6503
rect 4941 6447 5009 6503
rect 5065 6447 5133 6503
rect 5189 6447 5257 6503
rect 5313 6447 5381 6503
rect 5437 6447 5505 6503
rect 5561 6447 5629 6503
rect 5685 6447 5753 6503
rect 5809 6447 5877 6503
rect 5933 6447 6001 6503
rect 6057 6447 6125 6503
rect 6181 6447 6249 6503
rect 6305 6447 6373 6503
rect 6429 6447 6493 6503
rect 24 6379 6493 6447
rect 24 6323 4017 6379
rect 4073 6323 4141 6379
rect 4197 6323 4265 6379
rect 4321 6323 4389 6379
rect 4445 6323 4513 6379
rect 4569 6323 4637 6379
rect 4693 6323 4761 6379
rect 4817 6323 4885 6379
rect 4941 6323 5009 6379
rect 5065 6323 5133 6379
rect 5189 6323 5257 6379
rect 5313 6323 5381 6379
rect 5437 6323 5505 6379
rect 5561 6323 5629 6379
rect 5685 6323 5753 6379
rect 5809 6323 5877 6379
rect 5933 6323 6001 6379
rect 6057 6323 6125 6379
rect 6181 6323 6249 6379
rect 6305 6323 6373 6379
rect 6429 6323 6493 6379
rect 24 6255 6493 6323
rect 24 6199 4017 6255
rect 4073 6199 4141 6255
rect 4197 6199 4265 6255
rect 4321 6199 4389 6255
rect 4445 6199 4513 6255
rect 4569 6199 4637 6255
rect 4693 6199 4761 6255
rect 4817 6199 4885 6255
rect 4941 6199 5009 6255
rect 5065 6199 5133 6255
rect 5189 6199 5257 6255
rect 5313 6199 5381 6255
rect 5437 6199 5505 6255
rect 5561 6199 5629 6255
rect 5685 6199 5753 6255
rect 5809 6199 5877 6255
rect 5933 6199 6001 6255
rect 6057 6199 6125 6255
rect 6181 6199 6249 6255
rect 6305 6199 6373 6255
rect 6429 6199 6493 6255
rect 24 6131 6493 6199
rect 24 6075 4017 6131
rect 4073 6075 4141 6131
rect 4197 6075 4265 6131
rect 4321 6075 4389 6131
rect 4445 6075 4513 6131
rect 4569 6075 4637 6131
rect 4693 6075 4761 6131
rect 4817 6075 4885 6131
rect 4941 6075 5009 6131
rect 5065 6075 5133 6131
rect 5189 6075 5257 6131
rect 5313 6075 5381 6131
rect 5437 6075 5505 6131
rect 5561 6075 5629 6131
rect 5685 6075 5753 6131
rect 5809 6075 5877 6131
rect 5933 6075 6001 6131
rect 6057 6075 6125 6131
rect 6181 6075 6249 6131
rect 6305 6075 6373 6131
rect 6429 6075 6493 6131
rect 24 6007 6493 6075
rect 24 5951 4017 6007
rect 4073 5951 4141 6007
rect 4197 5951 4265 6007
rect 4321 5951 4389 6007
rect 4445 5951 4513 6007
rect 4569 5951 4637 6007
rect 4693 5951 4761 6007
rect 4817 5951 4885 6007
rect 4941 5951 5009 6007
rect 5065 5951 5133 6007
rect 5189 5951 5257 6007
rect 5313 5951 5381 6007
rect 5437 5951 5505 6007
rect 5561 5951 5629 6007
rect 5685 5951 5753 6007
rect 5809 5951 5877 6007
rect 5933 5951 6001 6007
rect 6057 5951 6125 6007
rect 6181 5951 6249 6007
rect 6305 5951 6373 6007
rect 6429 5951 6493 6007
rect 24 5884 6493 5951
rect 15454 6508 15826 6564
rect 15882 6508 15950 6564
rect 16006 6508 16074 6564
rect 16130 6508 16198 6564
rect 16254 6508 16322 6564
rect 16378 6508 16446 6564
rect 16502 6508 16570 6564
rect 16626 6508 16694 6564
rect 16750 6508 16818 6564
rect 16874 6508 17016 6564
rect 15454 6440 17016 6508
rect 15454 6384 15826 6440
rect 15882 6384 15950 6440
rect 16006 6384 16074 6440
rect 16130 6384 16198 6440
rect 16254 6384 16322 6440
rect 16378 6384 16446 6440
rect 16502 6384 16570 6440
rect 16626 6384 16694 6440
rect 16750 6384 16818 6440
rect 16874 6384 17016 6440
rect 15454 6316 17016 6384
rect 15454 6260 15826 6316
rect 15882 6260 15950 6316
rect 16006 6260 16074 6316
rect 16130 6260 16198 6316
rect 16254 6260 16322 6316
rect 16378 6260 16446 6316
rect 16502 6260 16570 6316
rect 16626 6260 16694 6316
rect 16750 6260 16818 6316
rect 16874 6260 17016 6316
rect 17284 7210 17907 7278
rect 17284 7154 17377 7210
rect 17433 7154 17501 7210
rect 17557 7154 17625 7210
rect 17681 7154 17749 7210
rect 17805 7154 17907 7210
rect 17284 7086 17907 7154
rect 17284 7030 17377 7086
rect 17433 7030 17501 7086
rect 17557 7030 17625 7086
rect 17681 7030 17749 7086
rect 17805 7030 17907 7086
rect 17284 6962 17907 7030
rect 17284 6906 17377 6962
rect 17433 6906 17501 6962
rect 17557 6906 17625 6962
rect 17681 6906 17749 6962
rect 17805 6906 17907 6962
rect 17284 6838 17907 6906
rect 17284 6782 17377 6838
rect 17433 6782 17501 6838
rect 17557 6782 17625 6838
rect 17681 6782 17749 6838
rect 17805 6782 17907 6838
rect 17284 6714 17907 6782
rect 17284 6658 17377 6714
rect 17433 6658 17501 6714
rect 17557 6658 17625 6714
rect 17681 6658 17749 6714
rect 17805 6658 17907 6714
rect 17284 6590 17907 6658
rect 17284 6534 17377 6590
rect 17433 6534 17501 6590
rect 17557 6534 17625 6590
rect 17681 6534 17749 6590
rect 17805 6534 17907 6590
rect 17284 6466 17907 6534
rect 17284 6410 17377 6466
rect 17433 6410 17501 6466
rect 17557 6410 17625 6466
rect 17681 6410 17749 6466
rect 17805 6410 17907 6466
rect 17284 6306 17907 6410
rect 15454 6192 17016 6260
rect 15454 6136 15826 6192
rect 15882 6136 15950 6192
rect 16006 6136 16074 6192
rect 16130 6136 16198 6192
rect 16254 6136 16322 6192
rect 16378 6136 16446 6192
rect 16502 6136 16570 6192
rect 16626 6136 16694 6192
rect 16750 6136 16818 6192
rect 16874 6136 17016 6192
rect 15454 6068 17016 6136
rect 15454 6012 15826 6068
rect 15882 6012 15950 6068
rect 16006 6012 16074 6068
rect 16130 6012 16198 6068
rect 16254 6012 16322 6068
rect 16378 6012 16446 6068
rect 16502 6012 16570 6068
rect 16626 6012 16694 6068
rect 16750 6012 16818 6068
rect 16874 6012 17016 6068
rect 15454 5944 17016 6012
rect 15454 5888 15826 5944
rect 15882 5888 15950 5944
rect 16006 5888 16074 5944
rect 16130 5888 16198 5944
rect 16254 5888 16322 5944
rect 16378 5888 16446 5944
rect 16502 5888 16570 5944
rect 16626 5888 16694 5944
rect 16750 5888 16818 5944
rect 16874 5888 17016 5944
rect 15454 5808 17016 5888
use std_buffer  std_buffer_0
timestamp 1765308861
transform 1 0 21358 0 -1 8992
box 1094 292 2782 3292
use reduction_mirror  X0
timestamp 1765308861
transform 1 0 -261 0 1 6308
box 261 -6308 25417 2408
use large_mimcap  X1
timestamp 1765308861
transform 1 0 11168 0 1 368
box -3514 -294 4286 7615
use schmitt_inverter  X2
timestamp 1765308861
transform 1 0 17635 0 1 8025
box 526 -2315 3059 685
use std_inverter  X3
timestamp 1765308861
transform 1 0 20638 0 -1 7361
box 265 -1350 1460 1650
<< labels >>
flabel metal5 s 803 8147 1003 8347 0 FreeSans 1600 0 0 0 VDD
port 1 nsew
flabel metal5 s 803 6188 1003 6388 0 FreeSans 1600 0 0 0 VSS
port 2 nsew
flabel metal2 s 24909 6342 25109 6542 0 FreeSans 1600 0 0 0 porb
port 3 nsew
flabel metal2 s 24908 6817 25108 7017 0 FreeSans 1600 0 0 0 por
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 25110 8710
string GDS_END 311492
string GDS_FILE ../gds/simple_por.gds.gz
string GDS_START 224738
<< end >>
