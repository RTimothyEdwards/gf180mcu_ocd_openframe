magic
tech gf180mcuD
magscale 1 10
timestamp 1765308861
<< metal1 >>
rect 1101 2992 1587 3292
rect 1249 2492 1384 2992
rect 1604 2862 1656 2883
rect 1604 2685 1656 2706
rect 1436 2599 1469 2651
rect 1521 2599 1554 2651
rect 1094 2163 1494 2185
rect 1094 2007 1316 2163
rect 1472 2007 1494 2163
rect 1094 1985 1494 2007
rect 1607 2159 1775 2167
rect 1607 2003 1613 2159
rect 1769 2003 1775 2159
rect 1607 1995 1775 2003
rect 2580 1980 2780 2180
rect 1222 592 1356 1483
rect 1424 1404 1524 1414
rect 1424 1352 1448 1404
rect 1500 1352 1524 1404
rect 1424 1342 1524 1352
rect 1553 1228 1605 1283
rect 1553 705 1605 760
rect 1111 292 1596 592
<< via1 >>
rect 1604 2706 1656 2862
rect 1469 2599 1521 2651
rect 1316 2007 1472 2163
rect 1613 2003 1769 2159
rect 1448 1352 1500 1404
rect 1553 760 1605 1228
<< metal2 >>
rect 1604 2885 1673 2888
rect 1602 2862 1673 2885
rect 1602 2706 1604 2862
rect 1656 2706 1673 2862
rect 1602 2683 1673 2706
rect 1446 2651 1544 2665
rect 1446 2599 1469 2651
rect 1521 2599 1544 2651
rect 1446 2584 1544 2599
rect 1446 2185 1513 2584
rect 1294 2163 1513 2185
rect 1604 2182 1673 2683
rect 1294 2007 1316 2163
rect 1472 2007 1513 2163
rect 1294 1985 1513 2007
rect 1435 1404 1513 1985
rect 1435 1352 1448 1404
rect 1500 1352 1513 1404
rect 1435 1327 1513 1352
rect 1578 2159 1788 2182
rect 1578 2003 1613 2159
rect 1769 2003 1788 2159
rect 1578 1982 1788 2003
rect 1578 1285 1649 1982
rect 1551 1228 1649 1285
rect 1551 760 1553 1228
rect 1605 760 1649 1228
rect 1551 703 1649 760
use std_inverter  X0
timestamp 1765308861
transform 1 0 1322 0 1 1642
box 265 -1350 1460 1650
use pmos_6p0_GUW2N9  XM2
timestamp 1765308861
transform 1 0 1474 0 1 1028
box -378 -586 368 586
use nmos_6p0_BUMBUS  XM3
timestamp 1765308861
transform 1 0 1505 0 1 2760
box -334 -332 334 332
<< labels >>
flabel metal1 s 1268 357 1468 557 0 FreeSans 1600 0 0 0 VDD
port 1 nsew
flabel metal1 s 1206 3043 1406 3243 0 FreeSans 1600 0 0 0 VSS
port 2 nsew
flabel metal1 s 1094 1985 1294 2185 0 FreeSans 1600 0 0 0 Vin
port 3 nsew
flabel metal1 s 2580 1980 2780 2180 0 FreeSans 1600 0 0 0 Vout
port 4 nsew
<< properties >>
string GDS_END 24024
string GDS_FILE ../gds/simple_por.gds.gz
string GDS_START 20646
<< end >>
