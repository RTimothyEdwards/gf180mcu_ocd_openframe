magic
tech gf180mcuD
magscale 1 10
timestamp 1765308861
<< error_p >>
rect -730 -255 -700 -209
rect -516 -255 -486 -209
rect -302 -255 -272 -209
rect -88 -255 -58 -209
rect 126 -255 156 -209
rect 340 -255 370 -209
rect 554 -255 584 -209
<< nwell >>
rect -1050 -486 980 486
<< hvpmos >>
rect -732 -176 -622 224
rect -518 -176 -408 224
rect -304 -176 -194 224
rect -90 -176 20 224
rect 124 -176 234 224
rect 338 -176 448 224
rect 552 -176 662 224
<< mvpdiff >>
rect -820 188 -732 224
rect -820 -140 -807 188
rect -761 -140 -732 188
rect -820 -176 -732 -140
rect -622 188 -518 224
rect -622 -140 -593 188
rect -547 -140 -518 188
rect -622 -176 -518 -140
rect -408 188 -304 224
rect -408 -140 -379 188
rect -333 -140 -304 188
rect -408 -176 -304 -140
rect -194 188 -90 224
rect -194 -140 -165 188
rect -119 -140 -90 188
rect -194 -176 -90 -140
rect 20 188 124 224
rect 20 -140 49 188
rect 95 -140 124 188
rect 20 -176 124 -140
rect 234 188 338 224
rect 234 -140 263 188
rect 309 -140 338 188
rect 234 -176 338 -140
rect 448 188 552 224
rect 448 -140 477 188
rect 523 -140 552 188
rect 448 -176 552 -140
rect 662 188 750 224
rect 662 -140 691 188
rect 737 -140 750 188
rect 662 -176 750 -140
<< mvpdiffc >>
rect -807 -140 -761 188
rect -593 -140 -547 188
rect -379 -140 -333 188
rect -165 -140 -119 188
rect 49 -140 95 188
rect 263 -140 309 188
rect 477 -140 523 188
rect 691 -140 737 188
<< mvnsubdiff >>
rect -964 387 894 400
rect -964 341 -810 387
rect 740 341 894 387
rect -964 328 894 341
rect -964 258 -892 328
rect -964 -258 -951 258
rect -905 -258 -892 258
rect 822 258 894 328
rect -964 -328 -892 -258
rect 822 -258 835 258
rect 881 -258 894 258
rect 822 -328 894 -258
rect -964 -400 894 -328
<< mvnsubdiffcont >>
rect -810 341 740 387
rect -951 -258 -905 258
rect 835 -258 881 258
<< polysilicon >>
rect -732 224 -622 268
rect -518 224 -408 268
rect -304 224 -194 268
rect -90 224 20 268
rect 124 224 234 268
rect 338 224 448 268
rect 552 224 662 268
rect -732 -209 -622 -176
rect -732 -255 -700 -209
rect -654 -255 -622 -209
rect -732 -268 -622 -255
rect -518 -209 -408 -176
rect -518 -255 -486 -209
rect -440 -255 -408 -209
rect -518 -268 -408 -255
rect -304 -209 -194 -176
rect -304 -255 -272 -209
rect -226 -255 -194 -209
rect -304 -268 -194 -255
rect -90 -209 20 -176
rect -90 -255 -58 -209
rect -12 -255 20 -209
rect -90 -268 20 -255
rect 124 -209 234 -176
rect 124 -255 156 -209
rect 202 -255 234 -209
rect 124 -268 234 -255
rect 338 -209 448 -176
rect 338 -255 370 -209
rect 416 -255 448 -209
rect 338 -268 448 -255
rect 552 -209 662 -176
rect 552 -255 584 -209
rect 630 -255 662 -209
rect 552 -268 662 -255
<< polycontact >>
rect -700 -255 -654 -209
rect -486 -255 -440 -209
rect -272 -255 -226 -209
rect -58 -255 -12 -209
rect 156 -255 202 -209
rect 370 -255 416 -209
rect 584 -255 630 -209
<< metal1 >>
rect -951 341 -810 387
rect 740 341 881 387
rect -951 258 -905 341
rect 835 258 881 341
rect -807 188 -761 222
rect -807 -174 -761 -140
rect -593 188 -547 222
rect -593 -174 -547 -140
rect -379 188 -333 222
rect -379 -174 -333 -140
rect -165 188 -119 222
rect -165 -174 -119 -140
rect 49 188 95 222
rect 49 -174 95 -140
rect 263 188 309 222
rect 263 -174 309 -140
rect 477 188 523 222
rect 477 -174 523 -140
rect 691 188 737 222
rect 691 -174 737 -140
rect -730 -255 -700 -209
rect -654 -255 -624 -209
rect -516 -255 -486 -209
rect -440 -255 -410 -209
rect -302 -255 -272 -209
rect -226 -255 -196 -209
rect -88 -255 -58 -209
rect -12 -255 18 -209
rect 126 -255 156 -209
rect 202 -255 232 -209
rect 340 -255 370 -209
rect 416 -255 446 -209
rect 554 -255 584 -209
rect 630 -255 660 -209
rect -951 -341 -905 -258
rect 835 -341 881 -258
rect -951 -387 881 -341
<< properties >>
string FIXED_BBOX -858 -364 858 364
string GDS_END 99246
string GDS_FILE ../gds/simple_por.gds.gz
string GDS_START 91946
<< end >>
