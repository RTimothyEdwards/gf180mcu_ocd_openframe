magic
tech gf180mcuD
magscale 1 10
timestamp 1764971740
<< checkpaint >>
rect -2001 2262 2303 2384
rect -2006 -1835 2303 2262
rect -2000 -1880 2303 -1835
rect -1951 -1885 2303 -1880
<< metal2 >>
rect 0 15194 59 15270
rect 222 15194 232 15270
rect 0 14673 59 14749
rect 222 14673 232 14749
rect 0 14444 59 14520
rect 222 14444 232 14520
rect 0 14302 59 14378
rect 222 14302 232 14378
rect 0 14160 59 14236
rect 222 14160 232 14236
rect 0 13800 59 13876
rect 222 13800 232 13876
rect 0 13589 59 13665
rect 222 13589 232 13665
rect 0 2132 59 2208
rect 222 2132 232 2208
rect 0 1986 59 2062
rect 222 1986 232 2062
rect 0 1840 59 1916
rect 222 1840 232 1916
rect 0 1694 59 1770
rect 222 1694 232 1770
rect 0 308 59 384
rect 222 308 232 384
rect 0 120 59 196
rect 222 120 232 196
<< via2 >>
rect 59 15194 222 15270
rect 59 14673 222 14749
rect 59 14444 222 14520
rect 59 14302 222 14378
rect 59 14160 222 14236
rect 59 13800 222 13876
rect 59 13589 222 13665
rect 59 2132 222 2208
rect 59 1986 222 2062
rect 59 1840 222 1916
rect 59 1694 222 1770
rect 59 308 222 384
rect 59 120 222 196
<< metal3 >>
rect 49 15194 59 15270
rect 222 15194 303 15270
rect 49 14673 59 14749
rect 222 14673 303 14749
rect 49 14444 59 14520
rect 222 14444 303 14520
rect 49 14302 59 14378
rect 222 14302 303 14378
rect 49 14160 59 14236
rect 222 14160 303 14236
rect 49 13800 59 13876
rect 222 13800 303 13876
rect 49 13589 59 13665
rect 222 13589 303 13665
rect 49 2132 59 2208
rect 222 2132 303 2208
rect 49 1986 59 2062
rect 222 1986 303 2062
rect 49 1840 59 1916
rect 222 1840 303 1916
rect 49 1694 59 1770
rect 222 1694 303 1770
rect 49 308 59 384
rect 222 308 303 384
rect 49 120 59 196
rect 222 120 303 196
<< properties >>
string flatten true
<< end >>
