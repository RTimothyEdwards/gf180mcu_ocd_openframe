magic
tech gf180mcuD
magscale 1 10
timestamp 1765305690
<< metal1 >>
rect 106424 103426 107485 103546
rect 90690 103110 92110 103122
rect 106426 103120 106546 103426
rect 90690 103010 90810 103110
rect 91140 103010 92110 103110
rect 90690 103002 92110 103010
rect 105317 103000 106546 103120
rect 106129 102642 107485 102762
rect 90690 102330 92110 102338
rect 106129 102336 106249 102642
rect 90690 102230 91270 102330
rect 91600 102230 92110 102330
rect 90690 102218 92110 102230
rect 105378 102216 106249 102336
rect 106424 101858 107485 101978
rect 90690 101540 92110 101554
rect 106426 101552 106546 101858
rect 90690 101440 90810 101540
rect 91140 101440 92110 101540
rect 90690 101434 92110 101440
rect 105378 101432 106546 101552
rect 106129 101074 107485 101194
rect 90690 100760 92110 100770
rect 106129 100768 106249 101074
rect 90690 100660 91270 100760
rect 91600 100660 92110 100760
rect 90690 100650 92110 100660
rect 105378 100648 106249 100768
rect 106424 100290 107485 100410
rect 90690 99980 92110 99986
rect 106426 99984 106546 100290
rect 90690 99880 90810 99980
rect 91140 99880 92110 99980
rect 90690 99866 92110 99880
rect 105378 99864 106546 99984
rect 106129 99506 107485 99626
rect 90690 99190 92110 99202
rect 106129 99200 106249 99506
rect 90690 99090 91270 99190
rect 91600 99090 92110 99190
rect 90690 99082 92110 99090
rect 105378 99080 106249 99200
rect 106424 98722 107485 98842
rect 90690 98410 92110 98418
rect 106426 98416 106546 98722
rect 90690 98310 90810 98410
rect 91140 98310 92110 98410
rect 90690 98298 92110 98310
rect 105378 98296 106546 98416
rect 106129 97938 107485 98058
rect 90690 97630 92110 97634
rect 106129 97632 106249 97938
rect 90690 97530 91270 97630
rect 91600 97530 92110 97630
rect 90690 97514 92110 97530
rect 105378 97512 106249 97632
rect 106424 97154 107485 97274
rect 90690 96840 92110 96850
rect 106426 96848 106546 97154
rect 90690 96740 90810 96840
rect 91140 96740 92110 96840
rect 90690 96730 92110 96740
rect 105378 96728 106546 96848
rect 106129 96370 107485 96490
rect 90690 96050 92110 96066
rect 106129 96064 106249 96370
rect 90690 95950 91270 96050
rect 91600 95950 92110 96050
rect 90690 95946 92110 95950
rect 105378 95944 106249 96064
rect 106424 95586 107485 95706
rect 90690 95270 92110 95282
rect 106426 95280 106546 95586
rect 90690 95170 90810 95270
rect 91140 95170 92110 95270
rect 90690 95162 92110 95170
rect 105378 95160 106546 95280
rect 106129 94802 107485 94922
rect 90690 94490 92110 94498
rect 106129 94496 106249 94802
rect 90690 94390 91270 94490
rect 91600 94390 92110 94490
rect 90690 94378 92110 94390
rect 105378 94376 106249 94496
rect 106424 94018 107485 94138
rect 90690 93700 92110 93714
rect 106426 93712 106546 94018
rect 90690 93600 90810 93700
rect 91140 93600 92110 93700
rect 90690 93594 92110 93600
rect 105378 93592 106546 93712
rect 106129 93234 107485 93354
rect 90690 92920 92110 92930
rect 106129 92928 106249 93234
rect 90690 92820 91270 92920
rect 91600 92820 92110 92920
rect 90690 92810 92110 92820
rect 105378 92808 106249 92928
rect 106424 92450 107485 92570
rect 90690 92140 92110 92146
rect 106426 92144 106546 92450
rect 90690 92040 90810 92140
rect 91140 92040 92110 92140
rect 90690 92026 92110 92040
rect 105379 92024 106546 92144
<< via1 >>
rect 90810 103010 91140 103110
rect 91270 102230 91600 102330
rect 90810 101440 91140 101540
rect 91270 100660 91600 100760
rect 90810 99880 91140 99980
rect 91270 99090 91600 99190
rect 90810 98310 91140 98410
rect 91270 97530 91600 97630
rect 90810 96740 91140 96840
rect 91270 95950 91600 96050
rect 90810 95170 91140 95270
rect 91270 94390 91600 94490
rect 90810 93600 91140 93700
rect 91270 92820 91600 92920
rect 90810 92040 91140 92140
<< metal2 >>
rect 90800 103110 91150 103220
rect 90800 103010 90810 103110
rect 91140 103010 91150 103110
rect 90800 101979 91150 103010
rect 90800 101540 91150 101859
rect 90800 101440 90810 101540
rect 91140 101440 91150 101540
rect 90800 100411 91150 101440
rect 90800 99980 91150 100291
rect 90800 99880 90810 99980
rect 91140 99880 91150 99980
rect 90800 98843 91150 99880
rect 90800 98410 91150 98723
rect 90800 98310 90810 98410
rect 91140 98310 91150 98410
rect 90800 97275 91150 98310
rect 90800 96840 91150 97155
rect 90800 96740 90810 96840
rect 91140 96740 91150 96840
rect 90800 95707 91150 96740
rect 90800 95270 91150 95587
rect 90800 95170 90810 95270
rect 91140 95170 91150 95270
rect 90800 94139 91150 95170
rect 90800 93700 91150 94019
rect 90800 93600 90810 93700
rect 91140 93600 91150 93700
rect 90800 92571 91150 93600
rect 90800 92140 91150 92451
rect 90800 92040 90810 92140
rect 91140 92040 91150 92140
rect 90800 91940 91150 92040
rect 91260 102775 91610 103220
rect 91260 102330 91610 102635
rect 91260 102230 91270 102330
rect 91600 102230 91610 102330
rect 91260 101207 91610 102230
rect 91260 100760 91610 101067
rect 91260 100660 91270 100760
rect 91600 100660 91610 100760
rect 91260 99639 91610 100660
rect 91260 99190 91610 99499
rect 91260 99090 91270 99190
rect 91600 99090 91610 99190
rect 91260 98071 91610 99090
rect 91260 97630 91610 97931
rect 91260 97530 91270 97630
rect 91600 97530 91610 97630
rect 91260 96503 91610 97530
rect 91260 96050 91610 96363
rect 91260 95950 91270 96050
rect 91600 95950 91610 96050
rect 91260 94935 91610 95950
rect 91260 94490 91610 94795
rect 91260 94390 91270 94490
rect 91600 94390 91610 94490
rect 91260 93367 91610 94390
rect 91260 92920 91610 93227
rect 91260 92820 91270 92920
rect 91600 92820 91610 92920
rect 91260 91940 91610 92820
<< via2 >>
rect 90800 101859 91150 101979
rect 90800 100291 91150 100411
rect 90800 98723 91150 98843
rect 90800 97155 91150 97275
rect 90800 95587 91150 95707
rect 90800 94019 91150 94139
rect 90800 92451 91150 92571
rect 91260 102635 91610 102775
rect 91260 101067 91610 101207
rect 91260 99499 91610 99639
rect 91260 97931 91610 98071
rect 91260 96363 91610 96503
rect 91260 94795 91610 94935
rect 91260 93227 91610 93367
<< metal3 >>
rect 88496 102635 91260 102775
rect 91610 102635 91640 102775
rect 88496 101859 90800 101979
rect 91150 101859 91170 101979
rect 88496 101067 91260 101207
rect 91610 101067 91640 101207
rect 88382 100291 90800 100411
rect 91150 100291 91170 100411
rect 88496 99499 91260 99639
rect 91610 99499 91640 99639
rect 88367 98723 90800 98843
rect 91150 98723 91170 98843
rect 88496 97931 91260 98071
rect 91610 97931 91640 98071
rect 88381 97155 90800 97275
rect 91150 97155 91170 97275
rect 88496 96363 91260 96503
rect 91610 96363 91640 96503
rect 88374 95587 90800 95707
rect 91150 95587 91170 95707
rect 88496 94795 91260 94935
rect 91610 94795 91640 94935
rect 88402 94019 90800 94139
rect 91150 94019 91170 94139
rect 88496 93227 91260 93367
rect 91610 93227 91640 93367
rect 88388 92451 90800 92571
rect 91150 92451 91170 92571
<< end >>
