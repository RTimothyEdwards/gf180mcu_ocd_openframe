* NGSPICE file created from caravel_openframe.ext - technology: gf180mcuD

.subckt POLY_SUB_FILL_1 a_597_223# a_685_131#
X0 a_685_131# a_597_223# cap_nmos_06v0 c_width=7u c_length=6u
X1 a_685_131# a_597_223# cap_nmos_06v0 c_width=7u c_length=6u
.ends

.subckt GF_NI_FILL10_1 VSS VDD DVSS DVDD
XPOLY_SUB_FILL_1_0[0] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[1] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[2] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[3] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[4] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[5] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[6] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[7] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[8] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[9] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[10] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[11] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[12] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[13] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[14] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[15] VSS VDD POLY_SUB_FILL_1
.ends

.subckt GF_NI_FILL10_0 DVSS DVDD VDD VSS
XGF_NI_FILL10_1_0 VSS VDD DVSS DVDD GF_NI_FILL10_1
.ends

.subckt gf180mcu_ocd_io__fill10 VDD VSS DVDD DVSS
XGF_NI_FILL10_0_0 DVSS DVDD VDD VSS GF_NI_FILL10_0
.ends

.subckt GF_NI_FILL10_1short VSS VDD DVSS DVDD
XPOLY_SUB_FILL_1_0[0] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[1] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[2] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[3] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[4] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[5] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[6] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[7] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[8] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[9] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[10] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[11] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[12] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[13] VSS VDD POLY_SUB_FILL_1
.ends

.subckt GF_NI_FILL10_0short DVSS DVDD VDD VSS
XGF_NI_FILL10_1_0 VSS VDD DVSS DVDD GF_NI_FILL10_1short
.ends

.subckt gf180mcu_as_sc_mcu7t3v3__decap_4 VDD VNW VPW VSS
X0 a_126_408# a_28_500# VSS VPW nfet_03v3 ad=0.44p pd=2.88u as=0.49p ps=2.98u w=1u l=1.03u
X1 VDD a_126_408# a_28_500# VNW pfet_03v3 ad=0.4752p pd=3.04u as=0.5292p ps=3.14u w=1.08u l=1.03u
.ends

.subckt gf180mcu_as_sc_mcu7t3v3__tiel_4 VDD VNW VPW VSS ZERO
X0 ZERO a_112_319# VSS VPW nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X1 a_112_319# a_112_319# VDD VNW pfet_03v3 ad=0.6072p pd=3.64u as=0.6072p ps=3.64u w=1.38u l=0.28u
.ends

.subckt gf180mcu_as_sc_mcu7t3v3__tieh_4 VDD VNW VPW VSS ONE
X0 a_112_319# a_112_319# VSS VPW nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X1 ONE a_112_319# VDD VNW pfet_03v3 ad=0.6072p pd=3.64u as=0.6072p ps=3.64u w=1.38u l=0.28u
.ends

.subckt gf180mcu_as_sc_mcu7t3v3__buff_12 VDD VNW VPW VSS A Y
X0 VSS a_172_68# Y VPW nfet_03v3 ad=0.985p pd=3.97u as=0.26p ps=1.52u w=1u l=0.28u
X1 VSS a_172_68# Y VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 VDD A a_172_68# VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X3 Y a_172_68# VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X4 Y a_172_68# VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X5 VDD a_172_68# Y VNW pfet_03v3 ad=1.3593p pd=4.73u as=0.3588p ps=1.9u w=1.38u l=0.28u
X6 a_172_68# A VSS VPW nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X7 VSS a_172_68# Y VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X8 VDD a_172_68# Y VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X9 Y a_172_68# VDD VNW pfet_03v3 ad=0.36915p pd=1.915u as=0.3588p ps=1.9u w=1.38u l=0.28u
X10 VDD a_172_68# Y VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X11 Y a_172_68# VSS VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X12 Y a_172_68# VSS VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X13 Y a_172_68# VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X14 Y a_172_68# VSS VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X15 a_172_68# A VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X16 VSS a_172_68# Y VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X17 VDD a_172_68# Y VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X18 VSS A a_172_68# VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X19 VSS a_172_68# Y VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X20 VSS a_172_68# Y VPW nfet_03v3 ad=0.26p pd=1.52u as=0.2675p ps=1.535u w=1u l=0.28u
X21 VDD A a_172_68# VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X22 Y a_172_68# VSS VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X23 Y a_172_68# VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X24 a_172_68# A VSS VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X25 Y a_172_68# VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X26 VDD a_172_68# Y VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X27 Y a_172_68# VSS VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X28 a_172_68# A VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.6072p ps=3.64u w=1.38u l=0.28u
X29 VDD a_172_68# Y VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.36915p ps=1.915u w=1.38u l=0.28u
X30 VSS A a_172_68# VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X31 Y a_172_68# VSS VPW nfet_03v3 ad=0.2675p pd=1.535u as=0.26p ps=1.52u w=1u l=0.28u
.ends

.subckt constant_block zero one vdd vss
Xgf180mcu_as_sc_mcu7t3v3__decap_4_0 vdd vdd vss vss gf180mcu_as_sc_mcu7t3v3__decap_4
Xgf180mcu_as_sc_mcu7t3v3__decap_4_1 vdd vdd vss vss gf180mcu_as_sc_mcu7t3v3__decap_4
Xgf180mcu_as_sc_mcu7t3v3__tiel_4_0 vdd vdd vss vss gf180mcu_as_sc_mcu7t3v3__buff_12_0/A
+ gf180mcu_as_sc_mcu7t3v3__tiel_4
Xgf180mcu_as_sc_mcu7t3v3__tieh_4_0 vdd vdd vss vss gf180mcu_as_sc_mcu7t3v3__buff_12_1/A
+ gf180mcu_as_sc_mcu7t3v3__tieh_4
Xgf180mcu_as_sc_mcu7t3v3__buff_12_1 vdd vdd vss vss gf180mcu_as_sc_mcu7t3v3__buff_12_1/A
+ one gf180mcu_as_sc_mcu7t3v3__buff_12
Xgf180mcu_as_sc_mcu7t3v3__buff_12_0 vdd vdd vss vss gf180mcu_as_sc_mcu7t3v3__buff_12_0/A
+ zero gf180mcu_as_sc_mcu7t3v3__buff_12
.ends

.subckt gf180mcu_ocd_io__fill10x VDD one zero DVDD DVSS VSS
XGF_NI_FILL10_0_0 DVSS DVDD VDD VSS GF_NI_FILL10_0short
Xconstant_block_0 zero one VDD VSS constant_block
.ends

.subckt lv_nand a_16960_50788# w_16870_51136# a_17113_51095# a_17024_51222# a_17252_51095#
X0 a_17204_50930# a_17113_51095# a_16960_50788# a_16960_50788# nfet_03v3 ad=0.114p pd=0.98u as=0.267p ps=2.09u w=0.6u l=0.28u
X1 a_17024_51222# a_17252_51095# a_17204_50930# a_16960_50788# nfet_03v3 ad=0.264p pd=2.08u as=0.114p ps=0.98u w=0.6u l=0.28u
X2 w_16870_51136# a_17113_51095# a_17024_51222# w_16870_51136# pfet_03v3 ad=0.333p pd=1.755u as=0.534p ps=3.29u w=1.2u l=0.28u
X3 a_17024_51222# a_17252_51095# w_16870_51136# w_16870_51136# pfet_03v3 ad=0.528p pd=3.28u as=0.333p ps=1.755u w=1.2u l=0.28u
.ends

.subckt pmos_6p0_esd_40 w_0_12# a_278_44# a_974_132# a_222_132#
X0 a_974_132# a_278_44# a_222_132# w_0_12# pfet_06v0_dss ad=0.1112n pd=85.56u as=11.2p ps=80.56u w=40u l=2.78u
.ends

.subckt comp018green_out_drv_pleg_4T_Y pmos_6p0_esd_40_0/w_0_12# pmos_6p0_esd_40_0/a_278_44#
+ pmos_6p0_esd_40_0/a_974_132# pmos_6p0_esd_40_0/a_222_132#
Xpmos_6p0_esd_40_0 pmos_6p0_esd_40_0/w_0_12# pmos_6p0_esd_40_0/a_278_44# pmos_6p0_esd_40_0/a_974_132#
+ pmos_6p0_esd_40_0/a_222_132# pmos_6p0_esd_40
.ends

.subckt comp018green_out_drv_pleg_4T_X pmos_6p0_esd_40_0/a_278_44# pmos_6p0_esd_40_1/w_0_12#
+ pmos_6p0_esd_40_0/a_222_132# pmos_6p0_esd_40_1/a_974_132# pmos_6p0_esd_40_1/a_278_44#
+ pmos_6p0_esd_40_1/a_222_132#
Xpmos_6p0_esd_40_0 pmos_6p0_esd_40_1/w_0_12# pmos_6p0_esd_40_0/a_278_44# pmos_6p0_esd_40_1/a_974_132#
+ pmos_6p0_esd_40_0/a_222_132# pmos_6p0_esd_40
Xpmos_6p0_esd_40_1 pmos_6p0_esd_40_1/w_0_12# pmos_6p0_esd_40_1/a_278_44# pmos_6p0_esd_40_1/a_974_132#
+ pmos_6p0_esd_40_1/a_222_132# pmos_6p0_esd_40
.ends

.subckt comp018green_out_paddrv_4T_PMOS_GROUP PMOS_4T_metal_stack_4/m1_340_0# a_2360_2800#
+ PMOS_4T_metal_stack_5/m1_340_0# a_4511_2800# PMOS_4T_metal_stack_5/m1_n44_0# PMOS_4T_metal_stack_1/m1_n44_0#
+ PMOS_4T_metal_stack_1/m1_340_0# PMOS_4T_metal_stack_2/m1_n44_0# a_9428_2800# a_7662_2800#
+ a_11201_2800# a_9815_2800# PMOS_4T_metal_stack_6/m1_340_0# PMOS_4T_metal_stack_2/m1_340_0#
+ PMOS_4T_metal_stack_3/m1_n44_0# a_6280_2800# a_2746_2800# a_974_2800# a_8049_2800#
+ a_5892_2800# PMOS_4T_metal_stack_3/m1_340_0# a_4120_2800# PMOS_4T_metal_stack_4/m1_n44_0#
+ w_n5_111#
Xcomp018green_out_drv_pleg_4T_Y_0 w_n5_111# a_4120_2800# PMOS_4T_metal_stack_1/m1_340_0#
+ PMOS_4T_metal_stack_2/m1_n44_0# comp018green_out_drv_pleg_4T_Y
Xcomp018green_out_drv_pleg_4T_Y_1 w_n5_111# a_9428_2800# PMOS_4T_metal_stack_4/m1_340_0#
+ PMOS_4T_metal_stack_5/m1_n44_0# comp018green_out_drv_pleg_4T_Y
Xcomp018green_out_drv_pleg_4T_Y_2 w_n5_111# a_2746_2800# PMOS_4T_metal_stack_1/m1_340_0#
+ PMOS_4T_metal_stack_1/m1_n44_0# comp018green_out_drv_pleg_4T_Y
Xcomp018green_out_drv_pleg_4T_Y_3 w_n5_111# a_8049_2800# PMOS_4T_metal_stack_4/m1_340_0#
+ PMOS_4T_metal_stack_4/m1_n44_0# comp018green_out_drv_pleg_4T_Y
Xcomp018green_out_drv_pleg_4T_X_0 a_4511_2800# w_n5_111# PMOS_4T_metal_stack_2/m1_n44_0#
+ PMOS_4T_metal_stack_2/m1_340_0# a_5892_2800# PMOS_4T_metal_stack_3/m1_n44_0# comp018green_out_drv_pleg_4T_X
Xcomp018green_out_drv_pleg_4T_X_1 a_9815_2800# w_n5_111# PMOS_4T_metal_stack_5/m1_n44_0#
+ PMOS_4T_metal_stack_5/m1_340_0# a_11201_2800# w_n5_111# comp018green_out_drv_pleg_4T_X
Xcomp018green_out_drv_pleg_4T_X_2 a_7662_2800# w_n5_111# PMOS_4T_metal_stack_4/m1_n44_0#
+ PMOS_4T_metal_stack_3/m1_340_0# a_6280_2800# PMOS_4T_metal_stack_3/m1_n44_0# comp018green_out_drv_pleg_4T_X
Xcomp018green_out_drv_pleg_4T_X_3 a_2360_2800# w_n5_111# PMOS_4T_metal_stack_1/m1_n44_0#
+ PMOS_4T_metal_stack_6/m1_340_0# a_974_2800# w_n5_111# comp018green_out_drv_pleg_4T_X
.ends

.subckt comp018green_out_drv_nleg_4T a_206_444# a_2080_444# a_2366_532# a_48_532#
+ a_436_532# VSUBS
X0 a_436_532# a_206_444# a_48_532# VSUBS nfet_06v0_dss ad=0.14364n pd=83.56u as=10.64p ps=76.56u w=38u l=3.78u
X1 a_2366_532# a_2080_444# a_436_532# VSUBS nfet_06v0_dss ad=10.64p pd=76.56u as=0.14364n ps=83.56u w=38u l=0.28u
.ends

.subckt comp018green_out_paddrv_4T_NMOS_GROUP GR_NMOS_4T_0/w_n1730_n583# a_7847_1028#
+ a_7373_1028# a_803_1028# nmos_4T_metal_stack_1/m1_n44_400# nmos_4T_metal_stack_2/m1_n44_400#
+ nmos_4T_metal_stack_3/m1_n44_400# nmos_4T_metal_stack_3/m1_430_401# a_2677_1028#
+ nmos_4T_metal_stack_1/m1_430_401# a_9721_1028# nmos_4T_metal_stack_2/m1_430_401#
+ nmos_4T_metal_stack_0/m1_n44_400# nmos_4T_metal_stack_4/m1_430_401# a_5499_1028#
+ a_3151_1028# VSUBS a_5025_1028# nmos_4T_metal_stack_4/m1_n44_400#
Xcomp018green_out_drv_nleg_4T_0 a_7847_1028# a_9721_1028# nmos_4T_metal_stack_0/m1_n44_400#
+ nmos_4T_metal_stack_3/m1_n44_400# nmos_4T_metal_stack_3/m1_430_401# VSUBS comp018green_out_drv_nleg_4T
Xcomp018green_out_drv_nleg_4T_1 a_5499_1028# a_7373_1028# nmos_4T_metal_stack_3/m1_n44_400#
+ nmos_4T_metal_stack_2/m1_n44_400# nmos_4T_metal_stack_2/m1_430_401# VSUBS comp018green_out_drv_nleg_4T
Xcomp018green_out_drv_nleg_4T_2 a_3151_1028# a_5025_1028# nmos_4T_metal_stack_2/m1_n44_400#
+ nmos_4T_metal_stack_1/m1_n44_400# nmos_4T_metal_stack_1/m1_430_401# VSUBS comp018green_out_drv_nleg_4T
Xcomp018green_out_drv_nleg_4T_3 a_803_1028# a_2677_1028# nmos_4T_metal_stack_1/m1_n44_400#
+ nmos_4T_metal_stack_4/m1_n44_400# nmos_4T_metal_stack_4/m1_430_401# VSUBS comp018green_out_drv_nleg_4T
.ends

.subckt comp018green_out_paddrv_16T comp018green_out_paddrv_4T_PMOS_GROUP_0/a_7662_2800#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/a_11201_2800# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_9428_2800#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_4/m1_n44_0# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_9815_2800#
+ m1_12305_8954# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_974_2800# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_6280_2800#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/a_2746_2800# m1_n360_8434# m1_1026_8954#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/w_n5_111# comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_1/m1_n44_0#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_5/m1_n44_0# m1_12305_9280#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/a_8049_2800# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_5892_2800#
+ comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_1/m1_n44_400# comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_2/m1_n44_400#
+ comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_3/m1_n44_400# m1_12305_9120#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/a_4120_2800# m1_1026_9280# comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_2/m1_n44_0#
+ m1_1026_9120# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_2360_2800# comp018green_out_paddrv_4T_NMOS_GROUP_0/VSUBS
+ m1_12305_9446# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_4511_2800# m2_1697_23319#
+ m1_1026_9446# comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_3/m1_n44_0#
Xcomp018green_out_paddrv_4T_PMOS_GROUP_0 m2_1697_23319# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_2360_2800#
+ m2_1697_23319# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_4511_2800# comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_5/m1_n44_0#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_1/m1_n44_0# m2_1697_23319#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_2/m1_n44_0# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_9428_2800#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/a_7662_2800# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_11201_2800#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/a_9815_2800# m2_1697_23319# m2_1697_23319#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_3/m1_n44_0# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_6280_2800#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/a_2746_2800# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_974_2800#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/a_8049_2800# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_5892_2800#
+ m2_1697_23319# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_4120_2800# comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_4/m1_n44_0#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/w_n5_111# comp018green_out_paddrv_4T_PMOS_GROUP
Xcomp018green_out_paddrv_4T_NMOS_GROUP_0 m1_n360_8434# m1_12305_9120# m1_12305_9280#
+ m1_1026_8954# comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_1/m1_n44_400#
+ comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_2/m1_n44_400# comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_3/m1_n44_400#
+ m2_1697_23319# m1_1026_9120# m2_1697_23319# m1_12305_8954# m2_1697_23319# comp018green_out_paddrv_4T_NMOS_GROUP_0/VSUBS
+ m2_1697_23319# m1_12305_9446# m1_1026_9280# comp018green_out_paddrv_4T_NMOS_GROUP_0/VSUBS
+ m1_1026_9446# comp018green_out_paddrv_4T_NMOS_GROUP_0/VSUBS comp018green_out_paddrv_4T_NMOS_GROUP
.ends

.subckt lvlshift_up a_18491_55181# a_18216_53410# a_18479_54386# a_18481_54667# w_18130_54691#
X0 w_18130_54691# a_18491_55181# a_18403_53764# w_18130_54691# pfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X1 a_18491_55181# a_18403_53764# w_18130_54691# w_18130_54691# pfet_06v0 ad=0.675p pd=3.9u as=0.39p ps=2.02u w=1.5u l=0.7u
X2 a_18216_53410# a_18479_54386# a_18403_53764# a_18216_53410# nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X3 a_18491_55181# a_18481_54667# a_18216_53410# a_18216_53410# nfet_06v0 ad=0.675p pd=3.9u as=0.39p ps=2.02u w=1.5u l=0.7u
.ends

.subckt comp018green_sigbuf_1 Z DVSS DVDD ZB lvlshift_up_0/a_18479_54386# lvlshift_up_0/a_18481_54667#
Xlvlshift_up_0 a_1605_310# DVSS lvlshift_up_0/a_18479_54386# lvlshift_up_0/a_18481_54667#
+ DVDD lvlshift_up
X0 DVSS Z ZB DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X1 Z a_1605_310# DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X2 ZB Z DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X3 DVDD Z ZB DVDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X4 ZB Z DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X5 DVDD a_1605_310# Z DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X6 Z a_1605_310# DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X7 DVSS a_1605_310# Z DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
.ends

.subckt comp018green_out_predrv SL SLB NDRIVE_X ENB DVSS A DVDD NDRIVE_Y PDRIVE_Y
+ PDRIVE_X EN
X0 a_1395_3267# ENB DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X1 DVDD a_1395_3267# PDRIVE_Y DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.7u
X2 NDRIVE_X a_335_226# DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.88u w=6u l=0.7u
X3 a_335_226# EN a_1395_3267# DVSS nfet_06v0 ad=2.64p pd=12.88u as=1.56p ps=6.52u w=6u l=0.7u
X4 NDRIVE_Y SL NDRIVE_X DVDD pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=12u l=0.7u
X5 DVSS a_335_226# NDRIVE_X DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X6 a_335_226# A DVDD DVDD pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=12u l=0.7u
X7 DVDD a_335_226# NDRIVE_Y DVDD pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=12u l=0.7u
X8 PDRIVE_X a_1395_3267# DVDD DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.7u
X9 PDRIVE_X DVDD PDRIVE_Y DVSS nfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X10 PDRIVE_Y SLB PDRIVE_X DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.88u w=6u l=0.7u
X11 NDRIVE_Y a_335_226# DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X12 PDRIVE_X SLB PDRIVE_Y DVSS nfet_06v0 ad=2.64p pd=12.88u as=1.56p ps=6.52u w=6u l=0.7u
X13 NDRIVE_Y a_335_226# DVDD DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.7u
X14 a_335_226# ENB a_1395_3267# DVDD pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=12u l=0.7u
X15 DVDD EN a_335_226# DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.7u
X16 NDRIVE_Y DVSS NDRIVE_X DVDD pfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X17 DVSS A a_1395_3267# DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.88u w=6u l=0.7u
X18 DVSS a_335_226# NDRIVE_Y DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X19 DVDD a_1395_3267# PDRIVE_X DVDD pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=12u l=0.7u
X20 PDRIVE_Y a_1395_3267# DVDD DVDD pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=12u l=0.7u
X21 PDRIVE_Y a_1395_3267# DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X22 DVSS a_1395_3267# PDRIVE_Y DVSS nfet_06v0 ad=2.64p pd=12.88u as=1.56p ps=6.52u w=6u l=0.7u
X23 NDRIVE_X SL NDRIVE_Y DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.7u
.ends

.subckt comp018green_out_sigbuf_a AB DVSS DVDD lvlshift_up_0/a_18479_54386# lvlshift_up_0/a_18481_54667#
Xlvlshift_up_0 a_1697_1072# DVSS lvlshift_up_0/a_18479_54386# lvlshift_up_0/a_18481_54667#
+ DVDD lvlshift_up
X0 AB a_1825_270# DVSS DVSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X1 AB a_1825_270# DVDD DVDD pfet_06v0 ad=2.64p pd=12.88u as=1.56p ps=6.52u w=6u l=0.7u
X2 DVSS a_1697_1072# a_1825_270# DVSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X3 DVDD a_1697_1072# a_1825_270# DVDD pfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.88u w=6u l=0.7u
.ends

.subckt comp018green_out_sigbuf_oe ENB DVDD DVSS EN lvlshift_up_0/a_18479_54386# lvlshift_up_0/a_18481_54667#
Xlvlshift_up_0 a_1783_1072# DVSS lvlshift_up_0/a_18479_54386# lvlshift_up_0/a_18481_54667#
+ DVDD lvlshift_up
X0 DVDD a_1783_1072# EN DVDD pfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.88u w=6u l=0.7u
X1 DVSS a_1783_1072# EN DVSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X2 ENB EN DVDD DVDD pfet_06v0 ad=2.64p pd=12.88u as=1.56p ps=6.52u w=6u l=0.7u
X3 ENB EN DVSS DVSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
.ends

.subckt lv_inv w_15980_51147# a_16280_50941# a_16119_51106# a_16066_50799#
X0 a_16280_50941# a_16119_51106# a_16066_50799# a_16066_50799# nfet_03v3 ad=0.264p pd=2.08u as=0.267p ps=2.09u w=0.6u l=0.28u
X1 a_16280_50941# a_16119_51106# w_15980_51147# w_15980_51147# pfet_03v3 ad=0.528p pd=3.28u as=0.558p ps=3.33u w=1.2u l=0.28u
.ends

.subckt comp018green_in_pupd A DVDD DVSS PU_B PD w_n83_53# a_506_484# a_6234_n7404#
X0 DVSS PD a_6278_n7492# DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X1 a_404_1044# a_7646_1324# w_n83_53# ppolyf_u r_width=0.8u r_length=35.7u
X2 a_404_2164# a_6278_n7492# w_n83_53# ppolyf_u r_width=0.8u r_length=35.7u
X3 DVDD a_6234_n7404# a_6278_n7492# DVDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X4 a_404_484# a_7646_764# w_n83_53# ppolyf_u r_width=0.8u r_length=35.7u
X5 a_404_1044# a_7646_764# w_n83_53# ppolyf_u r_width=0.8u r_length=35.7u
X6 a_404_2164# a_7646_1884# w_n83_53# ppolyf_u r_width=0.8u r_length=35.7u
X7 a_404_484# A w_n83_53# ppolyf_u r_width=0.8u r_length=23u
X8 a_404_1604# a_7646_1884# w_n83_53# ppolyf_u r_width=0.8u r_length=35.7u
X9 a_404_1604# a_7646_1324# w_n83_53# ppolyf_u r_width=0.8u r_length=35.7u
.ends

.subckt lv_passgate a_15637_45872# a_15397_45912# w_15280_46078# a_15366_45730# a_15492_45872#
+ a_15396_46108#
X0 a_15637_45872# a_15397_45912# a_15492_45872# a_15366_45730# nfet_03v3 ad=0.264p pd=2.08u as=0.267p ps=2.09u w=0.6u l=0.28u
X1 a_15637_45872# a_15396_46108# a_15492_45872# w_15280_46078# pfet_03v3 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.28u
.ends

.subckt comp018green_in_logic_pupd m1_1586_653# m1_1573_n494# m1_1324_578# m1_1842_n2708#
+ m1_1316_n577# a_1638_n204# w_1648_203# m1_1455_n1573#
Xlv_nand_4 a_1638_n204# w_1648_203# m1_1842_n2708# m1_1921_n496# m1_1909_n1494# lv_nand
Xlv_inv_0 w_1648_203# m1_1573_n494# m1_1921_n496# a_1638_n204# lv_inv
Xlv_inv_1 w_1648_203# m1_1586_653# m1_1910_652# a_1638_n204# lv_inv
Xlv_inv_2 w_1648_203# m1_1455_n1773# m1_1455_n1573# a_1638_n204# lv_inv
Xlv_passgate_0 m1_1909_n1494# m1_1455_n1573# w_1648_203# a_1638_n204# m1_1580_n1918#
+ m1_1455_n1773# lv_passgate
Xlv_inv_3 w_1648_203# m1_1580_n1918# m1_1842_n2708# a_1638_n204# lv_inv
Xlv_passgate_1 m1_1909_n1494# m1_1455_n1773# w_1648_203# a_1638_n204# m1_1842_n2708#
+ m1_1455_n1573# lv_passgate
Xlv_inv_5 w_1648_203# m1_1324_578# m1_1586_653# a_1638_n204# lv_inv
Xlv_inv_7 w_1648_203# m1_1316_n577# m1_1573_n494# a_1638_n204# lv_inv
Xlv_nand_0 a_1638_n204# w_1648_203# m1_1455_n1573# m1_1910_652# m1_1909_n1494# lv_nand
.ends

.subckt comp018green_sigbuf Z DVSS DVDD ZB IN INB
Xlvlshift_up_0 a_1561_310# DVSS IN INB DVDD lvlshift_up
X0 ZB Z DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X1 DVSS Z ZB DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X2 DVDD Z ZB DVDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X3 DVSS a_1561_310# Z DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X4 ZB Z DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X5 Z a_1561_310# DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X6 Z a_1561_310# DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X7 DVDD a_1561_310# Z DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
.ends

.subckt comp018green_in_drv DVDD A DVSS VDD VSS Z a_2771_580# a_1167_270# w_2679_1281#
+ a_923_1522# a_3067_747#
X0 VSS A a_n180_263# VSS nfet_06v0 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=0.7u
X1 a_n180_263# A VSS VSS nfet_06v0 ad=1.76p pd=8.88u as=1.04p ps=4.52u w=4u l=0.7u
X2 Z a_n180_263# a_1167_270# VSS nfet_06v0 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.7u
R0 VDD DVDD 0.000000
R1 VSS DVSS 0.000000
X3 a_1167_270# a_n180_263# Z VSS nfet_06v0 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.7u
X4 w_2679_1281# Z a_3067_747# w_2679_1281# pfet_03v3 ad=0.378p pd=1.94u as=0.378p ps=1.94u w=1.4u l=0.28u
X5 a_923_1522# a_n180_263# Z VDD pfet_06v0 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.7u
X6 a_2771_580# Z a_3067_747# a_2771_580# nfet_03v3 ad=0.162p pd=1.14u as=0.162p ps=1.14u w=0.6u l=0.28u
X7 a_3067_747# Z w_2679_1281# w_2679_1281# pfet_03v3 ad=0.378p pd=1.94u as=0.644p ps=3.72u w=1.4u l=0.28u
X8 a_3067_747# Z a_2771_580# a_2771_580# nfet_03v3 ad=0.162p pd=1.14u as=0.276p ps=2.12u w=0.6u l=0.28u
X9 a_3067_747# Z a_2771_580# a_2771_580# nfet_03v3 ad=0.162p pd=1.14u as=0.162p ps=1.14u w=0.6u l=0.28u
X10 a_3067_747# Z a_2771_580# a_2771_580# nfet_03v3 ad=0.162p pd=1.14u as=0.162p ps=1.14u w=0.6u l=0.28u
X11 a_2771_580# Z a_3067_747# a_2771_580# nfet_03v3 ad=0.276p pd=2.12u as=0.162p ps=1.14u w=0.6u l=0.28u
X12 a_2771_580# Z a_3067_747# a_2771_580# nfet_03v3 ad=0.162p pd=1.14u as=0.162p ps=1.14u w=0.6u l=0.28u
X13 Z a_n180_263# a_923_1522# VDD pfet_06v0 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.7u
X14 w_2679_1281# Z a_3067_747# w_2679_1281# pfet_03v3 ad=0.644p pd=3.72u as=0.378p ps=1.94u w=1.4u l=0.28u
X15 a_n180_263# A VDD VDD pfet_06v0 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.7u
X16 a_3067_747# Z w_2679_1281# w_2679_1281# pfet_03v3 ad=0.378p pd=1.94u as=0.378p ps=1.94u w=1.4u l=0.28u
X17 a_923_1522# a_n180_263# Z VDD pfet_06v0 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.7u
X18 w_2679_1281# Z a_3067_747# w_2679_1281# pfet_03v3 ad=0.378p pd=1.94u as=0.378p ps=1.94u w=1.4u l=0.28u
X19 a_3067_747# Z w_2679_1281# w_2679_1281# pfet_03v3 ad=0.378p pd=1.94u as=0.378p ps=1.94u w=1.4u l=0.28u
X20 Z a_n180_263# a_923_1522# VDD pfet_06v0 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.7u
.ends

.subckt comp018green_in_cms_smt IE CS DVDD A DVSS Z a_5355_608# m2_5364_1052#
X0 a_1887_280# IE DVSS DVSS nfet_06v0 ad=0.832p pd=3.72u as=0.832p ps=3.72u w=3.2u l=0.7u
X1 a_3115_338# a_1082_620# a_5355_608# DVSS nfet_06v0 ad=0.572p pd=3.48u as=0.572p ps=3.48u w=1.3u l=0.7u
X2 a_1082_620# a_599_280# Z DVDD pfet_06v0 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.7u
X3 DVSS CS a_599_280# DVSS nfet_06v0 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.7u
X4 DVSS a_1809_1797# a_3227_1730# DVDD pfet_06v0 ad=0.494p pd=2.42u as=0.836p ps=4.68u w=1.9u l=0.7u
X5 DVSS IE a_1887_280# DVSS nfet_06v0 ad=0.832p pd=3.72u as=0.832p ps=3.72u w=3.2u l=0.7u
X6 Z CS a_1809_1797# DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X7 Z IE DVDD DVDD pfet_06v0 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.7u
X8 Z a_599_280# a_1809_1797# DVDD pfet_06v0 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.7u
X9 a_1887_280# A a_3115_338# DVSS nfet_06v0 ad=0.689p pd=3.17u as=1.166p ps=6.18u w=2.65u l=0.7u
X10 DVDD CS a_1809_1797# DVDD pfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X11 a_3115_338# A a_1887_280# DVSS nfet_06v0 ad=0.689p pd=3.17u as=0.689p ps=3.17u w=2.65u l=0.7u
X12 Z A a_3227_1730# DVDD pfet_06v0 ad=0.559p pd=2.67u as=0.946p ps=5.18u w=2.15u l=0.7u
X13 a_3227_1730# A Z DVDD pfet_06v0 ad=0.946p pd=5.18u as=0.559p ps=2.67u w=2.15u l=0.7u
X14 DVSS a_599_280# a_1082_620# DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X15 a_1887_280# A a_3115_338# DVSS nfet_06v0 ad=0.689p pd=3.17u as=0.689p ps=3.17u w=2.65u l=0.7u
X16 DVDD A a_3227_1730# DVDD pfet_06v0 ad=0.494p pd=2.42u as=0.836p ps=4.68u w=1.9u l=0.7u
X17 a_1887_280# IE DVSS DVSS nfet_06v0 ad=1.408p pd=7.28u as=0.832p ps=3.72u w=3.2u l=0.7u
X18 Z A a_3115_338# DVSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X19 a_599_280# CS DVDD DVDD pfet_06v0 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=0.7u
X20 Z IE DVDD DVDD pfet_06v0 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.7u
X21 a_3115_338# A Z DVSS nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X22 DVDD IE Z DVDD pfet_06v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.7u
X23 a_3115_338# A a_1887_280# DVSS nfet_06v0 ad=1.166p pd=6.18u as=0.689p ps=3.17u w=2.65u l=0.7u
X24 a_1082_620# CS Z DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X25 a_3227_1730# A DVDD DVDD pfet_06v0 ad=0.836p pd=4.68u as=0.494p ps=2.42u w=1.9u l=0.7u
X26 a_3115_338# A Z DVSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X27 a_3227_1730# a_1809_1797# DVSS DVDD pfet_06v0 ad=0.836p pd=4.68u as=0.494p ps=2.42u w=1.9u l=0.7u
X28 a_599_280# CS DVSS DVSS nfet_06v0 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.7u
X29 DVDD CS a_599_280# DVDD pfet_06v0 ad=1.76p pd=8.88u as=1.04p ps=4.52u w=4u l=0.7u
X30 a_1887_280# IE DVSS DVSS nfet_06v0 ad=0.832p pd=3.72u as=1.408p ps=7.28u w=3.2u l=0.7u
X31 Z A a_3115_338# DVSS nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X32 a_1809_1797# CS DVDD DVDD pfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X33 DVSS IE a_1887_280# DVSS nfet_06v0 ad=0.832p pd=3.72u as=0.832p ps=3.72u w=3.2u l=0.7u
.ends

.subckt comp018green_inpath_cms_smt PAD CS PU comp018green_in_cms_smt_0/a_5355_608#
+ a_1390_1224# comp018green_in_logic_pupd_0/w_1648_203# comp018green_in_pupd_0/w_n83_53#
+ comp018green_in_pupd_0/A m3_9619_4882# m3_9619_3696# comp018green_in_pupd_0/DVSS
+ comp018green_in_pupd_0/DVDD comp018green_in_drv_0/VDD comp018green_in_drv_0/VSS
+ m1_12910_4326# VSUBS m1_10570_5335# comp018green_in_pupd_0/a_506_484# a_1390_2124#
+ w_n13_970# comp018green_sigbuf_3/DVSS comp018green_sigbuf_3/DVDD
Xlv_inv_14 w_n13_970# comp018green_sigbuf_1/IN a_1390_1224# VSUBS lv_inv
Xlv_inv_15 w_n13_970# comp018green_sigbuf_1/INB comp018green_sigbuf_1/IN VSUBS lv_inv
Xcomp018green_in_pupd_0 comp018green_in_pupd_0/A comp018green_in_pupd_0/DVDD comp018green_in_pupd_0/DVSS
+ comp018green_in_pupd_0/PU_B comp018green_sigbuf_0/ZB comp018green_in_pupd_0/w_n83_53#
+ comp018green_in_pupd_0/a_506_484# comp018green_sigbuf_2/Z comp018green_in_pupd
Xcomp018green_in_logic_pupd_0 comp018green_sigbuf_0/IN comp018green_sigbuf_2/IN comp018green_sigbuf_0/INB
+ PU comp018green_sigbuf_2/INB VSUBS comp018green_in_logic_pupd_0/w_1648_203# a_1390_2124#
+ comp018green_in_logic_pupd
Xcomp018green_sigbuf_0 comp018green_sigbuf_0/Z comp018green_sigbuf_3/DVSS comp018green_sigbuf_3/DVDD
+ comp018green_sigbuf_0/ZB comp018green_sigbuf_0/IN comp018green_sigbuf_0/INB comp018green_sigbuf
Xlv_inv_18 w_n13_970# comp018green_sigbuf_3/IN CS VSUBS lv_inv
Xlv_inv_19 w_n13_970# comp018green_sigbuf_3/INB comp018green_sigbuf_3/IN VSUBS lv_inv
Xcomp018green_sigbuf_1 comp018green_sigbuf_1/Z comp018green_sigbuf_3/DVSS comp018green_sigbuf_3/DVDD
+ comp018green_sigbuf_1/ZB comp018green_sigbuf_1/IN comp018green_sigbuf_1/INB comp018green_sigbuf
Xcomp018green_sigbuf_2 comp018green_sigbuf_2/Z comp018green_sigbuf_3/DVSS comp018green_sigbuf_3/DVDD
+ comp018green_sigbuf_2/ZB comp018green_sigbuf_2/IN comp018green_sigbuf_2/INB comp018green_sigbuf
Xcomp018green_sigbuf_3 comp018green_sigbuf_3/Z comp018green_sigbuf_3/DVSS comp018green_sigbuf_3/DVDD
+ comp018green_sigbuf_3/ZB comp018green_sigbuf_3/IN comp018green_sigbuf_3/INB comp018green_sigbuf
Xcomp018green_in_drv_0 comp018green_in_drv_0/VDD comp018green_in_drv_0/A comp018green_in_drv_0/VSS
+ comp018green_in_drv_0/VDD comp018green_in_drv_0/VSS comp018green_in_drv_0/Z VSUBS
+ VSUBS m1_10570_5335# m1_10570_5335# m1_12910_4326# comp018green_in_drv
Xcomp018green_in_cms_smt_0 comp018green_sigbuf_1/Z comp018green_sigbuf_3/Z comp018green_in_drv_0/VDD
+ PAD comp018green_in_drv_0/VSS comp018green_in_drv_0/A comp018green_in_cms_smt_0/a_5355_608#
+ PAD comp018green_in_cms_smt
D0 CS w_n13_970# diode_pd2nw_03v3 pj=4u area=1p
D1 a_1390_1224# w_n13_970# diode_pd2nw_03v3 pj=4u area=1p
D2 PU w_n13_970# diode_pd2nw_03v3 pj=4u area=1p
D3 a_1390_2124# w_n13_970# diode_pd2nw_03v3 pj=4u area=1p
.ends

.subckt comp018green_esd_cdm IP_IN PAD DVDD DVSS w_n86_n86# w_454_3720#
X0 PAD IP_IN DVDD ppolyf_u r_width=2.5u r_length=2.8u
D0 DVSS IP_IN diode_nd2ps_06v0 pj=42u area=20p
D1 IP_IN w_454_3720# diode_pd2nw_06v0 pj=42u area=20p
D2 DVSS IP_IN diode_nd2ps_06v0 pj=42u area=20p
X1 PAD IP_IN DVDD ppolyf_u r_width=2.5u r_length=2.8u
X2 PAD IP_IN DVDD ppolyf_u r_width=2.5u r_length=2.8u
X3 PAD IP_IN DVDD ppolyf_u r_width=2.5u r_length=2.8u
D3 IP_IN w_454_3720# diode_pd2nw_06v0 pj=42u area=20p
.ends

.subckt GF_NI_BI_T_BASE PD IE SL A OE CS PU PDRV0 PDRV1 Y ndrive_y_<0> ndrive_x_<0>
+ ndrive_x_<1> ndrive_Y_<1> ndrive_x_<2> ndrive_y_<2> ndrive_x_<3> ndrive_Y_<3> pdrive_x_<0>
+ pdrive_y_<0> pdrive_y_<1> pdrive_x_<1> pdrive_x_<2> pdrive_y_<2> pdrive_y_<3> pdrive_x_<3>
+ m3_1771_39126# w_11000_43887# comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_4/m1_n44_0#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/w_n5_111#
+ comp018green_inpath_cms_smt_0/m3_9619_4882# w_835_53274# comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_1/m1_n44_400#
+ comp018green_inpath_cms_smt_0/m3_9619_3696# comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_2/m1_n44_400#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_3/m1_n44_400#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_5/m1_n44_0#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_1/m1_n44_0#
+ comp018green_esd_cdm_0/w_454_3720# m3_10025_37504# PAD comp018green_inpath_cms_smt_0/comp018green_in_pupd_0/a_506_484#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_2/m1_n44_0#
+ a_12390_41548# m1_3608_46684# comp018green_esd_cdm_0/DVDD comp018green_inpath_cms_smt_0/comp018green_sigbuf_3/DVDD
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_3/m1_n44_0#
+ comp018green_sigbuf_1_0/VSUBS comp018green_esd_cdm_0/IP_IN comp018green_sigbuf_1_0/DVSS
+ comp018green_esd_cdm_0/DVSS comp018green_sigbuf_1_0/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VDD
+ a_882_55933# comp018green_inpath_cms_smt_0/m1_10570_5335# comp018green_inpath_cms_smt_0/VSUBS
+ w_11042_41027# comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/VSUBS
+ comp018green_out_predrv_3/DVDD w_13720_39292# comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS
Xlv_nand_2 comp018green_sigbuf_1_0/VSUBS w_13720_39292# OE m1_5236_36986# w_13720_39292#
+ lv_nand
Xlv_nand_3 comp018green_sigbuf_1_0/VSUBS w_13720_39292# OE m1_4812_38523# PDRV1 lv_nand
Xcomp018green_out_paddrv_16T_0 pdrive_x_<2> pdrive_x_<3> pdrive_y_<3> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_4/m1_n44_0#
+ pdrive_x_<3> ndrive_Y_<3> pdrive_x_<0> pdrive_x_<2> pdrive_y_<0> comp018green_out_predrv_3/DVDD
+ ndrive_x_<0> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/w_n5_111#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_1/m1_n44_0#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_5/m1_n44_0#
+ ndrive_y_<2> pdrive_y_<2> pdrive_x_<1> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_1/m1_n44_400#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_2/m1_n44_400#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_3/m1_n44_400#
+ ndrive_x_<3> pdrive_y_<1> ndrive_x_<1> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_2/m1_n44_0#
+ ndrive_y_<0> pdrive_x_<0> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/VSUBS
+ ndrive_x_<2> pdrive_x_<1> PAD ndrive_Y_<1> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_3/m1_n44_0#
+ comp018green_out_paddrv_16T
Xcomp018green_sigbuf_1_0 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/DVSS comp018green_sigbuf_1_0/DVDD
+ comp018green_sigbuf_1_0/ZB m1_9774_36986# m1_9537_37107# comp018green_sigbuf_1
Xcomp018green_out_predrv_0 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/ZB ndrive_x_<0>
+ comp018green_out_predrv_0/ENB comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_3/A
+ comp018green_out_predrv_3/DVDD ndrive_y_<0> pdrive_y_<0> pdrive_x_<0> comp018green_out_predrv_0/EN
+ comp018green_out_predrv
Xcomp018green_out_sigbuf_a_0 comp018green_out_predrv_3/A comp018green_sigbuf_1_0/DVSS
+ comp018green_sigbuf_1_0/DVDD m1_9178_38525# m1_9257_38818# comp018green_out_sigbuf_a
Xcomp018green_out_predrv_2 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/ZB ndrive_x_<2>
+ comp018green_out_predrv_3/ENB comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_3/A
+ comp018green_out_predrv_3/DVDD ndrive_y_<2> pdrive_y_<2> pdrive_x_<2> comp018green_out_predrv_3/EN
+ comp018green_out_predrv
Xcomp018green_out_predrv_1 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/ZB ndrive_x_<3>
+ comp018green_out_predrv_1/ENB comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_3/A
+ comp018green_out_predrv_3/DVDD ndrive_Y_<3> pdrive_y_<3> pdrive_x_<3> comp018green_out_predrv_1/EN
+ comp018green_out_predrv
Xcomp018green_out_sigbuf_oe_0 comp018green_out_predrv_0/ENB comp018green_sigbuf_1_0/DVDD
+ comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_0/EN m1_1184_38534# m1_1189_38806#
+ comp018green_out_sigbuf_oe
Xcomp018green_out_predrv_3 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/ZB ndrive_x_<1>
+ comp018green_out_predrv_3/ENB comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_3/A
+ comp018green_out_predrv_3/DVDD ndrive_Y_<1> pdrive_y_<1> pdrive_x_<1> comp018green_out_predrv_3/EN
+ comp018green_out_predrv
Xcomp018green_inpath_cms_smt_0 comp018green_esd_cdm_0/IP_IN CS PU comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VDD
+ IE w_11000_43887# m1_3608_46684# comp018green_esd_cdm_0/IP_IN comp018green_inpath_cms_smt_0/m3_9619_4882#
+ comp018green_inpath_cms_smt_0/m3_9619_3696# comp018green_esd_cdm_0/DVSS comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VDD
+ comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS
+ Y comp018green_inpath_cms_smt_0/VSUBS comp018green_inpath_cms_smt_0/m1_10570_5335#
+ comp018green_inpath_cms_smt_0/comp018green_in_pupd_0/a_506_484# PD w_835_53274#
+ comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS comp018green_inpath_cms_smt_0/comp018green_sigbuf_3/DVDD
+ comp018green_inpath_cms_smt
Xcomp018green_out_sigbuf_oe_2 comp018green_out_predrv_1/ENB comp018green_sigbuf_1_0/DVDD
+ comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_1/EN m1_5236_36986# m1_5084_37107#
+ comp018green_out_sigbuf_oe
Xcomp018green_out_sigbuf_oe_1 comp018green_out_predrv_3/ENB comp018green_sigbuf_1_0/DVDD
+ comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_3/EN m1_4812_38523# m1_4626_36747#
+ comp018green_out_sigbuf_oe
Xlv_inv_0 w_13720_39292# m1_1189_38806# m1_1184_38534# comp018green_sigbuf_1_0/VSUBS
+ lv_inv
Xlv_inv_1 w_13720_39292# m1_9257_38818# m1_9178_38525# comp018green_sigbuf_1_0/VSUBS
+ lv_inv
Xlv_inv_2 w_13720_39292# m1_9537_37107# m1_9774_36986# comp018green_sigbuf_1_0/VSUBS
+ lv_inv
Xlv_inv_3 w_13720_39292# m1_4626_36747# m1_4812_38523# comp018green_sigbuf_1_0/VSUBS
+ lv_inv
Xlv_inv_4 w_13720_39292# m1_9774_36986# SL comp018green_sigbuf_1_0/VSUBS lv_inv
Xlv_inv_6 w_13720_39292# m1_5084_37107# m1_5236_36986# comp018green_sigbuf_1_0/VSUBS
+ lv_inv
Xcomp018green_esd_cdm_0 comp018green_esd_cdm_0/IP_IN PAD comp018green_esd_cdm_0/DVDD
+ comp018green_esd_cdm_0/DVSS comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VDD
+ comp018green_esd_cdm_0/w_454_3720# comp018green_esd_cdm
Xlv_nand_0 comp018green_sigbuf_1_0/VSUBS w_13720_39292# OE m1_9178_38525# A lv_nand
Xlv_nand_1 comp018green_sigbuf_1_0/VSUBS w_13720_39292# OE m1_1184_38534# PDRV0 lv_nand
X0 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X1 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X2 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X3 a_882_55933# comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X4 a_882_55933# comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X5 a_12390_41548# comp018green_esd_cdm_0/DVSS cap_nmos_06v0 c_width=3u c_length=3u
X6 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X7 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X8 a_12390_41548# comp018green_esd_cdm_0/DVSS cap_nmos_06v0 c_width=3u c_length=3u
X9 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X10 a_12390_41548# comp018green_esd_cdm_0/DVSS cap_nmos_06v0 c_width=3u c_length=3u
X11 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
D0 comp018green_inpath_cms_smt_0/VSUBS OE diode_pd2nw_03v3 pj=1.92u area=0.2304p
D1 comp018green_inpath_cms_smt_0/VSUBS OE diode_pd2nw_03v3 pj=1.92u area=0.2304p
D2 comp018green_inpath_cms_smt_0/VSUBS OE diode_pd2nw_03v3 pj=1.92u area=0.2304p
D3 comp018green_inpath_cms_smt_0/VSUBS w_11000_43887# diode_pd2nw_03v3 pj=1.92u area=0.2304p
D4 A w_11042_41027# diode_pd2nw_03v3 pj=4u area=1p
D5 SL w_11042_41027# diode_pd2nw_03v3 pj=4u area=1p
X12 a_12390_41548# comp018green_esd_cdm_0/DVSS cap_nmos_06v0 c_width=3u c_length=3u
D6 comp018green_inpath_cms_smt_0/VSUBS PDRV0 diode_pd2nw_03v3 pj=1.92u area=0.2304p
D7 comp018green_inpath_cms_smt_0/VSUBS PDRV1 diode_pd2nw_03v3 pj=1.92u area=0.2304p
X13 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
.ends

.subckt gf180mcu_ocd_io__bi_a DVDD PDRV0 PDRV1 PU VDD ANA A IE PAD SL Y OE PD CS VSS
+ DVSS
XGF_NI_BI_T_BASE_0 PD IE SL A OE CS PU PDRV0 PDRV1 Y GF_NI_BI_T_BASE_0/ndrive_y_<0>
+ GF_NI_BI_T_BASE_0/ndrive_x_<0> GF_NI_BI_T_BASE_0/ndrive_x_<1> GF_NI_BI_T_BASE_0/ndrive_Y_<1>
+ GF_NI_BI_T_BASE_0/ndrive_x_<2> GF_NI_BI_T_BASE_0/ndrive_y_<2> GF_NI_BI_T_BASE_0/ndrive_x_<3>
+ GF_NI_BI_T_BASE_0/ndrive_Y_<3> GF_NI_BI_T_BASE_0/pdrive_x_<0> GF_NI_BI_T_BASE_0/pdrive_y_<0>
+ GF_NI_BI_T_BASE_0/pdrive_y_<1> GF_NI_BI_T_BASE_0/pdrive_x_<1> GF_NI_BI_T_BASE_0/pdrive_x_<2>
+ GF_NI_BI_T_BASE_0/pdrive_y_<2> GF_NI_BI_T_BASE_0/pdrive_y_<3> GF_NI_BI_T_BASE_0/pdrive_x_<3>
+ VDD VDD DVDD DVDD VDD VDD DVSS VSS DVSS DVSS DVDD DVDD DVDD VSS PAD a_3151_58293#
+ DVDD DVDD DVDD DVDD DVDD DVDD VSS ANA DVSS DVSS DVDD DVDD DVDD VDD VSS VDD DVSS
+ DVDD VDD DVSS GF_NI_BI_T_BASE
.ends

.subckt POLY_SUB_FILL a_1165_n91# a_1077_1#
X0 a_1165_n91# a_1077_1# cap_nmos_06v0 c_width=1.5u c_length=1.5u
X1 a_1165_n91# a_1077_1# cap_nmos_06v0 c_width=1.5u c_length=1.5u
.ends

.subckt GF_NI_FILL5_1 VSS VDD DVSS DVDD
XPOLY_SUB_FILL_0[0] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[1] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[2] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[3] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[4] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[5] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[6] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[7] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[8] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[9] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[10] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[11] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[12] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[13] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[14] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[15] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[16] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[17] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[18] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[19] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[20] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[21] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[22] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[23] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[24] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[25] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[26] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[27] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[28] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[29] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[30] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[31] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[32] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[33] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[34] VDD VSS POLY_SUB_FILL
.ends

.subckt GF_NI_FILL5_0 DVSS DVDD VDD VSS
XGF_NI_FILL5_1_0 VSS VDD DVSS DVDD GF_NI_FILL5_1
.ends

.subckt gf180mcu_ocd_io__fill5 VDD VSS DVDD DVSS
XGF_NI_FILL5_0_0 DVSS DVDD VDD VSS GF_NI_FILL5_0
.ends

.subckt comp018green_esd_rc_v5p0 VRC VPLUS VMINUS
X0 a_353_2269# a_13226_1989# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X1 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X2 a_353_3389# a_13226_3109# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X3 a_353_2829# a_13226_3109# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X4 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X5 a_353_1709# a_13226_1989# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X6 a_353_1709# a_13226_1429# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X7 a_353_2829# a_13226_2549# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X8 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X9 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X10 VRC a_13226_3669# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X11 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X12 a_353_1149# a_13226_1429# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X13 VPLUS a_13226_869# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X14 a_353_2269# a_13226_2549# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X15 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X16 a_353_3389# a_13226_3669# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X17 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X18 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X19 a_353_1149# a_13226_869# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
.ends

.subckt nmos_clamp_20_50_4_DVDD a_582_632# w_n51_n51# a_1237_1481#
X0 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X1 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X2 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X3 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X4 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X5 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X6 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X7 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X8 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X9 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X10 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X11 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X12 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X13 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X14 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X15 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X16 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X17 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X18 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X19 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X20 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X21 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X22 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X23 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X24 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X25 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X26 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X27 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X28 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X29 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X30 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X31 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X32 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X33 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X34 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X35 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X36 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X37 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X38 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X39 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X40 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X41 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X42 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X43 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X44 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
X45 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X46 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X47 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X48 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X49 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X50 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X51 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X52 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X53 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X54 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
X55 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
X56 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X57 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X58 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X59 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X60 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X61 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X62 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X63 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X64 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X65 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X66 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X67 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X68 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X69 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X70 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X71 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X72 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X73 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X74 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X75 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X76 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X77 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X78 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X79 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
.ends

.subckt comp018green_esd_clamp_v5p0_DVDD comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VMINUS
Xcomp018green_esd_rc_v5p0_0 comp018green_esd_rc_v5p0_0/VRC comp018green_esd_rc_v5p0_0/VPLUS
+ comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0
Xnmos_clamp_20_50_4_DVDD_0 comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VPLUS
+ a_4685_27917# nmos_clamp_20_50_4_DVDD
X0 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X1 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X2 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X3 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X4 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X5 a_3781_27917# a_2805_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X6 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.7u
X7 comp018green_esd_rc_v5p0_0/VMINUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X8 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X9 a_3781_27917# a_2805_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.7u
X10 comp018green_esd_rc_v5p0_0/VMINUS a_2805_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X11 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X12 a_3781_27917# a_2805_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X13 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X14 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X15 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X16 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X17 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X18 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X19 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X20 comp018green_esd_rc_v5p0_0/VMINUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X21 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X22 comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VRC a_2805_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X23 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X24 a_2805_27917# comp018green_esd_rc_v5p0_0/VRC comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=2.2p pd=10.88u as=2.2p ps=10.88u w=5u l=0.7u
X25 comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VRC a_2805_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X26 comp018green_esd_rc_v5p0_0/VMINUS a_2805_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X27 a_2805_27917# comp018green_esd_rc_v5p0_0/VRC comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.7u
X28 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X29 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X30 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X31 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X32 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.7u
X33 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X34 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X35 a_3781_27917# a_2805_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.7u
X36 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X37 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X38 comp018green_esd_rc_v5p0_0/VMINUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.7u
X39 a_2805_27917# comp018green_esd_rc_v5p0_0/VRC comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X40 a_3781_27917# a_2805_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X41 comp018green_esd_rc_v5p0_0/VMINUS a_2805_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X42 comp018green_esd_rc_v5p0_0/VPLUS a_2805_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X43 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
.ends

.subckt GF_NI_VDD_BASE DVSS DVDD VSS m3_9927_12842# m3_7265_56043# m3_5168_14436#
+ m3_7265_52842# m3_12297_33636# m3_2798_11242# m3_12297_56043# m3_2798_17636# m3_9927_1636#
+ m3_12297_52842# m3_7265_8036# m3_12861_28842# m3_9927_33636# m3_7265_4836# m3_7874_28842#
+ m3_12861_24036# m3_12861_54442# m3_10244_14436# m3_4851_27242# m3_9927_56043# m3_5168_11242#
+ m3_9927_52842# m3_7874_24036# m3_7874_54442# m3_2798_30436# m3_12861_20836# m3_12861_43242#
+ m3_5168_17636# m3_12861_41642# m3_7265_48042# m3_2481_27242# m3_7874_20836# m3_9927_8036#
+ m3_7874_43242# m3_12297_1636# m3_7874_41642# m3_4851_12842# m3_7265_44842# m3_9927_4836#
+ m3_12297_48042# m3_10244_11242# m3_5168_30436# m3_2481_12842# m3_12297_44842# m3_10244_17636#
+ m3_2481_1636# m3_2798_28842# m3_9927_48042# m3_4851_33636# m3_12297_8036# m3_12861_14436#
+ m3_2798_24036# m3_2798_54442# m3_4851_56043# m3_9927_44842# m3_12297_4836# m3_4851_52842#
+ m3_7874_14436# m3_2481_33636# m3_10244_30436# m3_2798_20836# m3_2798_43242# m3_2798_41642#
+ m3_4851_1636# m3_2481_56043# m3_5168_28842# m3_2481_8036# m3_2481_52842# m3_7265_27242#
+ m3_5168_24036# m3_2481_4836# m3_5168_54442# m3_12861_11242# m3_5168_20836# m3_5168_43242#
+ m3_12297_27242# m3_12861_17636# m3_7874_11242# m3_5168_41642# m3_4851_8036# m3_10244_28842#
+ m3_4851_48042# m3_7265_12842# m3_7874_17636# m3_4851_4836# m3_10244_24036# m3_2798_14436#
+ m3_10244_54442# m3_4851_44842# m3_9927_27242# m3_12297_12842# m3_2481_48042# VDD
+ m3_12861_30436# m3_10244_20836# m3_10244_43242# m3_7265_1636# m3_10244_41642# m3_2481_44842#
+ m3_7874_30436# m3_7265_33636#
Xcomp018green_esd_clamp_v5p0_DVDD_0 VDD VSS comp018green_esd_clamp_v5p0_DVDD
D0 VSS VDD diode_nd2ps_06v0 pj=82u area=40p
X0 VDD VSS cap_nmos_06v0 c_width=15u c_length=15u
D1 VSS VDD diode_nd2ps_06v0 pj=82u area=40p
D2 VSS VDD diode_nd2ps_06v0 pj=82u area=40p
D3 VSS VDD diode_nd2ps_06v0 pj=82u area=40p
X1 VDD VSS cap_nmos_06v0 c_width=15u c_length=15u
X2 VDD VSS cap_nmos_06v0 c_width=15u c_length=15u
X3 VDD VSS cap_nmos_06v0 c_width=15u c_length=15u
.ends

.subckt gf180mcu_ocd_io__vdd DVDD DVSS VDD VSS
XGF_NI_VDD_BASE_0 DVSS DVDD VSS DVSS DVSS DVDD DVSS DVSS DVDD DVSS DVDD DVSS DVSS
+ DVSS DVDD DVSS DVSS DVDD DVDD DVDD DVDD DVSS DVSS DVDD DVSS DVDD DVDD DVDD DVDD
+ DVDD DVDD DVDD DVSS DVSS DVDD DVSS DVDD DVSS DVDD DVSS DVSS DVSS DVSS DVDD DVDD
+ DVSS DVSS DVDD DVSS DVDD DVSS DVSS DVSS DVDD DVDD DVDD DVSS DVSS DVSS DVSS DVDD
+ DVSS DVDD DVDD DVDD DVDD DVSS DVSS DVDD DVSS DVSS DVSS DVDD DVSS DVDD DVDD DVDD
+ DVDD DVSS DVDD DVDD DVDD DVSS DVDD DVSS DVSS DVDD DVSS DVDD DVDD DVDD DVSS DVSS
+ DVSS DVSS VDD DVDD DVDD DVDD DVSS DVDD DVSS DVDD DVSS GF_NI_VDD_BASE
.ends

.subckt pmos_6p0_GUW2N9 a_50_n324# w_n378_n586# a_n148_n324# a_n60_n368#
X0 a_50_n324# a_n60_n368# a_n148_n324# w_n378_n586# pfet_05v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.55u
.ends

.subckt nmos_6p0_BUMBUS a_n302_n300# a_n70_n168# a_n158_n76# a_70_n76#
X0 a_70_n76# a_n70_n168# a_n158_n76# a_n302_n300# nfet_05v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt pmos_6p0_MUW2NR a_n52_n524# w_n480_n786# a_162_n524# a_n162_n568# a_n250_n524#
+ a_52_n568#
X0 a_n52_n524# a_n162_n568# a_n250_n524# w_n480_n786# pfet_05v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.55u
X1 a_162_n524# a_52_n568# a_n52_n524# w_n480_n786# pfet_05v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.55u
.ends

.subckt nmos_6p0_BUMBJU a_n158_n276# a_n302_n500# a_n70_n368# a_70_n276#
X0 a_70_n276# a_n70_n368# a_n158_n276# a_n302_n500# nfet_05v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
.ends

.subckt std_inverter VDD Vin Vout VSS
XXM0 Vout VDD VDD Vin VDD Vin pmos_6p0_MUW2NR
XXM1 VSS VSS Vin Vout nmos_6p0_BUMBJU
.ends

.subckt std_buffer VDD Vin Vout VSS
XXM2 X0/Vin VDD VDD Vin pmos_6p0_GUW2N9
XXM3 VSS Vin VSS X0/Vin nmos_6p0_BUMBUS
XX0 VDD X0/Vin Vout VSS std_inverter
.ends

.subckt nmos_6p0_BJPB5U a_n70_n268# a_n158_n224# a_70_n224# a_n302_n400#
X0 a_70_n224# a_n70_n268# a_n158_n224# a_n302_n400# nfet_05v0 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.7u
.ends

.subckt pmos_6p0_EYEQQM a_n304_n268# a_n622_n176# a_234_n176# a_n408_n176# a_124_n268#
+ a_n732_n268# w_n1050_n486# a_n518_n268# a_n90_n268# a_662_n176# a_n820_n176# a_448_n176#
+ a_n194_n176# a_552_n268# a_20_n176# a_338_n268#
X0 a_448_n176# a_338_n268# a_234_n176# w_n1050_n486# pfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.55u
X1 a_n194_n176# a_n304_n268# a_n408_n176# w_n1050_n486# pfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.55u
X2 a_n408_n176# a_n518_n268# a_n622_n176# w_n1050_n486# pfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.55u
X3 a_662_n176# a_552_n268# a_448_n176# w_n1050_n486# pfet_05v0 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.55u
X4 a_20_n176# a_n90_n268# a_n194_n176# w_n1050_n486# pfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.55u
X5 a_n622_n176# a_n732_n268# a_n820_n176# w_n1050_n486# pfet_05v0 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.55u
X6 a_234_n176# a_124_n268# a_20_n176# w_n1050_n486# pfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.55u
.ends

.subckt nmos_6p0_B4TB5U a_n70_n268# a_70_n176# a_n158_n176# a_n302_n400#
X0 a_70_n176# a_n70_n268# a_n158_n176# a_n302_n400# nfet_05v0 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.7u
.ends

.subckt pmos_6p0_CYEQN4 a_n138_n176# a_60_n176# a_n50_n268# w_n368_n486#
X0 a_60_n176# a_n50_n268# a_n138_n176# w_n368_n486# pfet_05v0 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.55u
.ends

.subckt nmos_6p0_BJXXPT a_662_n268# a_n314_n268# a_n70_n268# a_n418_n224# a_n1034_n400#
+ a_n174_n224# a_802_n224# a_n802_n268# a_n890_n224# a_n662_n224# a_418_n268# a_174_n268#
+ a_558_n224# a_314_n224# a_70_n224# a_n558_n268#
X0 a_n662_n224# a_n802_n268# a_n890_n224# a_n1034_n400# nfet_05v0 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.7u
X1 a_n174_n224# a_n314_n268# a_n418_n224# a_n1034_n400# nfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.7u
X2 a_802_n224# a_662_n268# a_558_n224# a_n1034_n400# nfet_05v0 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.7u
X3 a_n418_n224# a_n558_n268# a_n662_n224# a_n1034_n400# nfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.7u
X4 a_70_n224# a_n70_n268# a_n174_n224# a_n1034_n400# nfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.7u
X5 a_314_n224# a_174_n268# a_70_n224# a_n1034_n400# nfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.7u
X6 a_558_n224# a_418_n268# a_314_n224# a_n1034_n400# nfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.7u
.ends

.subckt ppolyf_u_1k_6p0_TRTT7C a_7600_n2622# a_5360_2500# a_2560_n2622# a_3120_n2622#
+ a_n5280_2500# a_8720_n2622# a_4800_2500# a_12080_n2622# a_3680_n2622# a_n8080_n2622#
+ a_600_2500# a_4240_n2622# a_n4720_2500# a_9840_n2622# a_6200_2500# a_5640_2500#
+ a_n1640_n2622# a_n10040_n2622# a_5360_n2622# a_n6120_2500# a_11800_n2622# a_880_2500#
+ a_n2200_n2622# a_n5560_2500# a_n240_2500# a_n7800_n2622# a_n240_n2622# a_n2760_n2622#
+ a_n11160_n2622# a_6480_n2622# a_7040_2500# a_6480_2500# a_n3320_n2622# a_7040_n2622#
+ a_n8920_n2622# a_n3880_n2622# a_n12280_n2622# a_5920_2500# a_n4440_n2622# a_8160_n2622#
+ a_n6400_2500# a_n5840_2500# a_n520_2500# a_n5000_n2622# a_1160_2500# a_7320_2500#
+ a_n5560_n2622# a_6760_2500# a_9280_n2622# a_320_n2622# a_n1080_2500# a_10120_n2622#
+ a_1720_n2622# a_n6120_n2622# a_n7240_2500# a_880_n2622# a_n1080_n2622# a_n6680_2500#
+ a_10680_n2622# a_n6680_n2622# a_8160_2500# a_11240_n2622# a_2840_n2622# a_n7240_n2622#
+ a_2000_2500# a_n800_2500# a_3400_n2622# a_1440_2500# a_n8080_2500# a_7600_2500#
+ a_n1360_2500# a_n8360_n2622# a_3960_n2622# a_4520_n2622# a_n7520_2500# a_n6960_2500#
+ a_2280_2500# a_n9480_n2622# a_n10040_2500# a_9000_2500# a_8440_2500# a_5640_n2622#
+ a_n1920_n2622# a_n10320_n2622# a_7880_2500# a_10120_2500# a_6200_n2622# a_1720_2500#
+ a_n8360_2500# a_n10880_n2622# a_n520_n2622# a_n2200_2500# a_1160_n2622# a_n1640_2500#
+ a_n11440_n2622# a_6760_n2622# a_9280_2500# a_n3600_n2622# a_n7800_2500# a_n12000_n2622#
+ a_7320_n2622# a_3120_2500# a_n10320_2500# a_2560_2500# a_2280_n2622# a_7880_n2622#
+ a_n3040_2500# a_8720_2500# a_n2480_2500# a_n4720_n2622# a_8440_n2622# a_10400_2500#
+ a_n9200_2500# a_n12492_n2834# a_n8640_2500# a_40_n2622# a_9000_n2622# a_n1920_2500#
+ a_n11160_2500# a_n5840_n2622# a_9560_n2622# a_9560_2500# a_10400_n2622# a_600_n2622#
+ a_11240_2500# a_n6400_n2622# a_3400_2500# a_10680_2500# a_n9480_2500# a_n10600_2500#
+ a_10960_n2622# a_2840_2500# a_n1360_n2622# a_5080_n2622# a_n3320_2500# a_n6960_n2622#
+ a_11520_n2622# a_n2760_2500# a_n7520_n2622# a_n8920_2500# a_12080_2500# a_n2480_n2622#
+ a_n12000_2500# a_4240_2500# a_3680_2500# a_n11440_2500# a_n3040_n2622# a_n10880_2500#
+ a_n4160_2500# a_n8640_n2622# a_9840_2500# a_11520_2500# a_4800_n2622# a_10960_2500#
+ a_n9200_n2622# a_n9760_2500# a_n4160_n2622# a_5080_2500# a_40_2500# a_n3600_2500#
+ a_n9760_n2622# a_n12280_2500# a_n10600_n2622# a_5920_n2622# a_n5280_n2622# a_4520_2500#
+ a_3960_2500# a_n5000_2500# a_n11720_2500# a_1440_n2622# a_320_2500# a_n800_n2622#
+ a_n4440_2500# a_n11720_n2622# a_n3880_2500# a_11800_2500# a_2000_n2622#
X0 a_n6400_2500# a_n6400_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X1 a_n3320_2500# a_n3320_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X2 a_1720_2500# a_1720_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X3 a_7040_2500# a_7040_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X4 a_n5840_2500# a_n5840_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X5 a_9560_2500# a_9560_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X6 a_n10040_2500# a_n10040_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X7 a_5080_2500# a_5080_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X8 a_n3880_2500# a_n3880_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X9 a_n1360_2500# a_n1360_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X10 a_2000_2500# a_2000_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X11 a_4520_2500# a_4520_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X12 a_n10600_2500# a_n10600_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X13 a_n9200_2500# a_n9200_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X14 a_n6120_2500# a_n6120_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X15 a_11520_2500# a_11520_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X16 a_12080_2500# a_12080_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X17 a_n8640_2500# a_n8640_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X18 a_n4160_2500# a_n4160_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X19 a_2560_2500# a_2560_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X20 a_n6680_2500# a_n6680_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X21 a_7320_2500# a_7320_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X22 a_9840_2500# a_9840_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X23 a_n10320_2500# a_n10320_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X24 a_n2200_2500# a_n2200_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X25 a_5360_2500# a_5360_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X26 a_n1640_2500# a_n1640_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X27 a_4800_2500# a_4800_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X28 a_7880_2500# a_7880_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X29 a_n10880_2500# a_n10880_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X30 a_n9480_2500# a_n9480_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X31 a_n8920_2500# a_n8920_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X32 a_11800_2500# a_11800_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X33 a_2840_2500# a_2840_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X34 a_n4440_2500# a_n4440_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X35 a_8160_2500# a_8160_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X36 a_n11160_2500# a_n11160_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X37 a_n6960_2500# a_n6960_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X38 a_320_2500# a_320_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X39 a_7600_2500# a_7600_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X40 a_n5000_2500# a_n5000_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X41 a_n2480_2500# a_n2480_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X42 a_n1920_2500# a_n1920_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X43 a_3120_2500# a_3120_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X44 a_5640_2500# a_5640_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X45 a_n9760_2500# a_n9760_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X46 a_n7240_2500# a_n7240_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X47 a_880_2500# a_880_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X48 a_10120_2500# a_10120_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X49 a_1160_2500# a_1160_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X50 a_3680_2500# a_3680_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X51 a_n5280_2500# a_n5280_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X52 a_n240_2500# a_n240_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X53 a_40_2500# a_40_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X54 a_n7800_2500# a_n7800_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X55 a_n4720_2500# a_n4720_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X56 a_8440_2500# a_8440_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X57 a_10680_2500# a_10680_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X58 a_n11440_2500# a_n11440_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X59 a_600_2500# a_600_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X60 a_n2760_2500# a_n2760_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X61 a_n800_2500# a_n800_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X62 a_3400_2500# a_3400_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X63 a_6480_2500# a_6480_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X64 a_n8080_2500# a_n8080_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X65 a_5920_2500# a_5920_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X66 a_n12000_2500# a_n12000_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X67 a_n7520_2500# a_n7520_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X68 a_10400_2500# a_10400_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X69 a_1440_2500# a_1440_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X70 a_3960_2500# a_3960_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X71 a_n5560_2500# a_n5560_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X72 a_n3040_2500# a_n3040_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X73 a_n520_2500# a_n520_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X74 a_6200_2500# a_6200_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X75 a_9280_2500# a_9280_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X76 a_10960_2500# a_10960_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X77 a_n12280_2500# a_n12280_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X78 a_8720_2500# a_8720_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X79 a_n11720_2500# a_n11720_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X80 a_n3600_2500# a_n3600_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X81 a_n1080_2500# a_n1080_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X82 a_4240_2500# a_4240_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X83 a_6760_2500# a_6760_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X84 a_n8360_2500# a_n8360_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X85 a_9000_2500# a_9000_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X86 a_11240_2500# a_11240_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
X87 a_2280_2500# a_2280_n2622# a_n12492_n2834# ppolyf_u_1k_6p0 r_width=1u r_length=25u
.ends

.subckt pmos_6p0_HUEQQM a_375_n176# a_265_n268# a_n810_n268# a_n596_n268# a_803_n176#
+ a_n272_n176# a_589_n176# a_161_n176# a_693_n268# a_n58_n176# a_479_n268# a_51_n268#
+ a_n382_n268# w_n1128_n486# a_n168_n268# a_n898_n176# a_n700_n176# a_n486_n176#
X0 a_375_n176# a_265_n268# a_161_n176# w_n1128_n486# pfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.55u
X1 a_n272_n176# a_n382_n268# a_n486_n176# w_n1128_n486# pfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.55u
X2 a_n700_n176# a_n810_n268# a_n898_n176# w_n1128_n486# pfet_05v0 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.55u
X3 a_589_n176# a_479_n268# a_375_n176# w_n1128_n486# pfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.55u
X4 a_n486_n176# a_n596_n268# a_n700_n176# w_n1128_n486# pfet_05v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.55u
X5 a_161_n176# a_51_n268# a_n58_n176# w_n1128_n486# pfet_05v0 ad=0.52p pd=2.52u as=0.545p ps=2.545u w=2u l=0.55u
X6 a_n58_n176# a_n168_n268# a_n272_n176# w_n1128_n486# pfet_05v0 ad=0.545p pd=2.545u as=0.52p ps=2.52u w=2u l=0.55u
X7 a_803_n176# a_693_n268# a_589_n176# w_n1128_n486# pfet_05v0 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.55u
.ends

.subckt reduction_mirror VDD Vout VSS
Xnmos_6p0_BJPB5U_0 m2_1393_n86# VSS m2_3858_n195# VSS nmos_6p0_BJPB5U
Xpmos_6p0_EYEQQM_0 m2_4433_1027# VDD VDD m2_4433_1027# m2_4433_1027# m2_4433_1027#
+ VDD m2_4433_1027# m2_4433_1027# VDD m2_4433_1027# m2_4433_1027# VDD m2_4433_1027#
+ m2_4433_1027# m2_4433_1027# pmos_6p0_EYEQQM
XXM0 m1_2517_n836# VSS m2_607_119# VSS nmos_6p0_B4TB5U
XXM1 m2_3432_1017# m2_1393_n86# m2_607_119# VDD pmos_6p0_CYEQN4
Xpmos_6p0_CYEQN4_0 m2_6726_1023# Vout m2_3858_n195# VDD pmos_6p0_CYEQN4
XXM3 m2_607_119# m2_921_1004# m2_607_119# VDD pmos_6p0_CYEQN4
XXM4 VDD m2_3432_1017# m2_921_1004# VDD pmos_6p0_CYEQN4
XXM7 VDD m2_6726_1023# m2_4433_1027# VDD pmos_6p0_CYEQN4
XXM9 m2_3858_n195# m2_4433_1027# m2_3858_n195# VDD pmos_6p0_CYEQN4
Xnmos_6p0_BJXXPT_0 m2_1393_n86# m2_1393_n86# m2_1393_n86# m2_1393_n86# VSS VSS VSS
+ m2_1393_n86# m2_1393_n86# VSS m2_1393_n86# m2_1393_n86# m2_1393_n86# VSS m2_1393_n86#
+ m2_1393_n86# nmos_6p0_BJXXPT
Xppolyf_u_1k_6p0_TRTT7C_0 m1_20155_n6001# m1_18197_n836# m1_15115_n6001# m1_15675_n6001#
+ m1_7557_n836# m1_21275_n6001# m1_17637_n836# m1_24635_n6001# m1_16235_n6001# m1_4475_n6001#
+ m1_13157_n836# m1_16795_n6001# m1_8117_n836# m1_22395_n6001# m1_18757_n836# m1_18197_n836#
+ m1_11195_n6001# m1_2795_n6001# m1_17915_n6001# m1_6437_n836# m1_24635_n6001# m1_13717_n836#
+ m1_10635_n6001# m1_6997_n836# m1_12597_n836# m1_5035_n6001# m1_12315_n6001# m1_10075_n6001#
+ m1_1675_n6001# m1_19035_n6001# m1_19877_n836# m1_19317_n836# m1_9515_n6001# m1_19595_n6001#
+ m1_3915_n6001# m1_8955_n6001# m1_555_n6001# m1_18757_n836# m1_8395_n6001# m1_20715_n6001#
+ m1_6437_n836# m1_6997_n836# m1_12037_n836# m1_7835_n6001# m1_13717_n836# m1_19877_n836#
+ m1_7275_n6001# m1_19317_n836# m1_21835_n6001# m1_12875_n6001# m1_11477_n836# m1_22955_n6001#
+ m1_14555_n6001# m1_6715_n6001# m1_5317_n836# m1_13435_n6001# m1_11755_n6001# m1_5877_n836#
+ m1_23515_n6001# m1_6155_n6001# m1_20997_n836# m1_24075_n6001# m1_15675_n6001# m1_5595_n6001#
+ m1_14837_n836# m1_12037_n836# m1_16235_n6001# m1_14277_n836# m1_4757_n836# m1_20437_n836#
+ m1_11477_n836# m1_4475_n6001# m1_16795_n6001# m1_17355_n6001# m1_5317_n836# m1_5877_n836#
+ m1_14837_n836# m1_3355_n6001# m1_2517_n836# m1_21557_n836# m1_20997_n836# m1_18475_n6001#
+ m1_10635_n6001# m1_2235_n6001# m1_20437_n836# m1_22677_n836# m1_19035_n6001# m1_14277_n836#
+ m1_4197_n836# m1_1675_n6001# m1_12315_n6001# m1_10357_n836# m1_13995_n6001# m1_10917_n836#
+ m1_1115_n6001# m1_19595_n6001# m1_22117_n836# m1_8955_n6001# m1_4757_n836# m1_555_n6001#
+ m1_20155_n6001# m1_15957_n836# m1_2517_n836# m1_15397_n836# m1_15115_n6001# m1_20715_n6001#
+ m1_9797_n836# m1_21557_n836# m1_10357_n836# m1_7835_n6001# m1_21275_n6001# m1_23237_n836#
+ m1_3637_n836# VSS m1_4197_n836# m1_12875_n6001# m1_21835_n6001# m1_10917_n836# m1_1397_n836#
+ m1_6715_n6001# m1_22395_n6001# m1_22117_n836# m1_22955_n6001# m1_13435_n6001# m1_23797_n836#
+ m1_6155_n6001# m1_15957_n836# m1_23237_n836# m1_3077_n836# m1_1957_n836# m1_23515_n6001#
+ m1_15397_n836# m1_11195_n6001# m1_17915_n6001# m1_9237_n836# m1_5595_n6001# m1_24075_n6001#
+ m1_9797_n836# m1_5035_n6001# m1_3637_n836# VDD m1_10075_n6001# m1_837_n836# m1_17077_n836#
+ m1_16517_n836# m1_1397_n836# m1_9515_n6001# m1_1957_n836# m1_8677_n836# m1_3915_n6001#
+ m1_22677_n836# m1_24357_n836# m1_17355_n6001# m1_23797_n836# m1_3355_n6001# m1_3077_n836#
+ m1_8395_n6001# m1_17637_n836# m1_12597_n836# m1_9237_n836# m1_2795_n6001# VSS m1_2235_n6001#
+ m1_18475_n6001# m1_7275_n6001# m1_17077_n836# m1_16517_n836# m1_7557_n836# m1_837_n836#
+ m1_13995_n6001# m1_13157_n836# m1_11755_n6001# m1_8117_n836# m1_1115_n6001# m1_8677_n836#
+ m1_24357_n836# m1_14555_n6001# ppolyf_u_1k_6p0_TRTT7C
Xpmos_6p0_HUEQQM_0 m2_921_1004# m2_921_1004# m2_921_1004# m2_921_1004# m2_921_1004#
+ VDD VDD VDD m2_921_1004# m2_921_1004# m2_921_1004# m2_921_1004# m2_921_1004# VDD
+ m2_921_1004# m2_921_1004# VDD m2_921_1004# pmos_6p0_HUEQQM
.ends

.subckt mim_2p0fF_8KW78G m4_n1220_n1120# m4_n1100_n1000#
X0 m4_n1100_n1000# m4_n1220_n1120# cap_mim_2f0_m4m5_noshield c_width=10u c_length=10u
.ends

.subckt large_mimcap In VSS
XXC1[0|0] VSS In mim_2p0fF_8KW78G
XXC1[1|0] VSS In mim_2p0fF_8KW78G
XXC1[2|0] VSS In mim_2p0fF_8KW78G
XXC1[0|1] VSS In mim_2p0fF_8KW78G
XXC1[1|1] VSS In mim_2p0fF_8KW78G
XXC1[2|1] VSS In mim_2p0fF_8KW78G
XXC1[0|2] VSS In mim_2p0fF_8KW78G
XXC1[1|2] VSS In mim_2p0fF_8KW78G
XXC1[2|2] VSS In mim_2p0fF_8KW78G
.ends

.subckt pmos_6p0_UXEQNM a_n60_n168# a_n148_n76# w_n378_n386# a_50_n76#
X0 a_50_n76# a_n60_n168# a_n148_n76# w_n378_n386# pfet_05v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
.ends

.subckt nmos_6p0_L3YBEV a_n188_n724# a_100_n724# a_n332_n900# a_n100_n768#
X0 a_100_n724# a_n100_n768# a_n188_n724# a_n332_n900# nfet_05v0 ad=3.08p pd=14.88u as=3.08p ps=14.88u w=7u l=1u
.ends

.subckt pmos_6p0_9YEQN4 a_50_n576# w_n378_n886# a_n148_n576# a_n60_n668#
X0 a_50_n576# a_n60_n668# a_n148_n576# w_n378_n886# pfet_05v0 ad=2.64p pd=12.88u as=2.64p ps=12.88u w=6u l=0.55u
.ends

.subckt pmos_6p0_9859UL a_n288_n26# a_n200_n118# a_200_n26# w_n518_n336#
X0 a_200_n26# a_n200_n118# a_n288_n26# w_n518_n336# pfet_05v0 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=2u
.ends

.subckt schmitt_inverter VDD VSS Vin Vout
Xpmos_6p0_UXEQNM_0 Vin m1_1072_n872# VDD Vout pmos_6p0_UXEQNM
XX6 m1_1243_n1927# VDD VSS Vout nmos_6p0_L3YBEV
Xnmos_6p0_BJPB5U_0 Vin m1_1243_n1927# Vout VSS nmos_6p0_BJPB5U
XXM1 m1_1072_n872# VDD VDD Vin pmos_6p0_9YEQN4
XXM3 Vin VSS m1_1243_n1927# VSS nmos_6p0_BJPB5U
XXM5 m1_1072_n872# Vout VSS VDD pmos_6p0_9859UL
.ends

.subckt simple_por VDD porb por VSS
Xstd_buffer_0 VDD X3/Vin por VSS std_buffer
XX0 VDD X1/In VSS reduction_mirror
XX1 X1/In VSS large_mimcap
XX2 VDD VSS X1/In X3/Vin schmitt_inverter
XX3 VDD X3/Vin porb VSS std_inverter
.ends

.subckt nmos_clamp_20_50_4_DVSS a_582_632# w_n51_n51# a_1237_1481#
X0 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X1 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X2 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X3 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X4 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X5 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X6 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X7 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X8 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X9 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X10 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X11 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X12 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X13 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X14 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X15 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X16 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X17 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X18 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X19 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X20 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X21 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X22 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X23 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X24 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X25 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X26 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X27 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X28 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X29 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X30 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X31 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X32 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X33 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X34 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X35 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X36 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X37 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X38 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X39 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X40 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X41 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X42 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X43 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X44 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
X45 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X46 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X47 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X48 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X49 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X50 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X51 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X52 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X53 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X54 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
X55 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
X56 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X57 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X58 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X59 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X60 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X61 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X62 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X63 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X64 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X65 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X66 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X67 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X68 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X69 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X70 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X71 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X72 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X73 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X74 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X75 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X76 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X77 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X78 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X79 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
.ends

.subckt comp018green_esd_clamp_v5p0_DVSS comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VMINUS
Xcomp018green_esd_rc_v5p0_0 comp018green_esd_rc_v5p0_0/VRC comp018green_esd_rc_v5p0_0/VPLUS
+ comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0
Xnmos_clamp_20_50_4_DVSS_0 comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VPLUS
+ a_4685_27917# nmos_clamp_20_50_4_DVSS
X0 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X1 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X2 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X3 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X4 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X5 a_3781_27917# a_2805_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X6 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.7u
X7 comp018green_esd_rc_v5p0_0/VMINUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X8 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X9 a_3781_27917# a_2805_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.7u
X10 comp018green_esd_rc_v5p0_0/VMINUS a_2805_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X11 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X12 a_3781_27917# a_2805_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X13 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X14 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X15 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X16 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X17 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X18 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X19 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X20 comp018green_esd_rc_v5p0_0/VMINUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X21 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X22 comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VRC a_2805_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X23 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X24 a_2805_27917# comp018green_esd_rc_v5p0_0/VRC comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=2.2p pd=10.88u as=2.2p ps=10.88u w=5u l=0.7u
X25 comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VRC a_2805_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X26 comp018green_esd_rc_v5p0_0/VMINUS a_2805_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X27 a_2805_27917# comp018green_esd_rc_v5p0_0/VRC comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.7u
X28 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X29 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X30 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X31 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X32 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.7u
X33 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X34 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X35 a_3781_27917# a_2805_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.7u
X36 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X37 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X38 comp018green_esd_rc_v5p0_0/VMINUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.7u
X39 a_2805_27917# comp018green_esd_rc_v5p0_0/VRC comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X40 a_3781_27917# a_2805_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X41 comp018green_esd_rc_v5p0_0/VMINUS a_2805_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X42 comp018green_esd_rc_v5p0_0/VPLUS a_2805_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X43 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
.ends

.subckt GF_NI_DVSS_BASE DVDD m2_2292_38400# a_12742_47643# DVSS comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS
Xcomp018green_esd_clamp_v5p0_DVSS_0 comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS
+ DVSS comp018green_esd_clamp_v5p0_DVSS
D0 DVSS comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS diode_nd2ps_06v0 pj=82u area=40p
X0 comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS DVSS cap_nmos_06v0 c_width=15u c_length=15u
D1 DVSS comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS diode_nd2ps_06v0 pj=82u area=40p
D2 DVSS comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS diode_nd2ps_06v0 pj=82u area=40p
D3 DVSS comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS diode_nd2ps_06v0 pj=82u area=40p
X1 comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS DVSS cap_nmos_06v0 c_width=15u c_length=15u
X2 comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS DVSS cap_nmos_06v0 c_width=15u c_length=15u
X3 comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS DVSS cap_nmos_06v0 c_width=15u c_length=15u
.ends

.subckt gf180mcu_ocd_io__dvss DVDD DVSS VDD VSS
XGF_NI_DVSS_BASE_0 DVDD VDD VSS DVSS DVDD GF_NI_DVSS_BASE
.ends

.subckt GF_NI_DVDD_BASE DVSS a_246_47643# a_13001_27179# m2_2279_36800# comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0/VMINUS
+ DVDD
Xcomp018green_esd_clamp_v5p0_DVDD_0 DVDD comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0/VMINUS
+ comp018green_esd_clamp_v5p0_DVDD
D0 comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0/VMINUS DVDD diode_nd2ps_06v0 pj=82u area=40p
X0 DVDD comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0/VMINUS cap_nmos_06v0 c_width=15u c_length=15u
D1 comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0/VMINUS DVDD diode_nd2ps_06v0 pj=82u area=40p
D2 comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0/VMINUS DVDD diode_nd2ps_06v0 pj=82u area=40p
D3 comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0/VMINUS DVDD diode_nd2ps_06v0 pj=82u area=40p
X1 DVDD comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0/VMINUS cap_nmos_06v0 c_width=15u c_length=15u
X2 DVDD comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0/VMINUS cap_nmos_06v0 c_width=15u c_length=15u
X3 DVDD comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0/VMINUS cap_nmos_06v0 c_width=15u c_length=15u
.ends

.subckt gf180mcu_ocd_io__dvdd VDD VSS DVDD DVSS
XGF_NI_DVDD_BASE_0 DVSS VSS VSS VSS DVSS DVDD GF_NI_DVDD_BASE
.ends

.subckt moscap_corner_1 a_5519_6541# a_5519_529# a_4904_32#
X0 a_5519_529# a_4904_32# cap_nmos_06v0 c_width=25u c_length=10u
X1 a_5519_6541# a_4904_32# cap_nmos_06v0 c_width=25u c_length=10u
X2 a_5519_529# a_4904_32# cap_nmos_06v0 c_width=25u c_length=10u
X3 a_5519_6541# a_4904_32# cap_nmos_06v0 c_width=25u c_length=10u
.ends

.subckt moscap_corner VMINUS a_647_6541# a_647_529#
X0 a_647_6541# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X1 a_647_529# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X2 a_647_6541# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X3 a_647_529# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X4 a_647_529# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X5 a_647_6541# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X6 a_647_6541# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X7 a_647_529# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
.ends

.subckt nmos_clamp_20_50_4 a_582_632# w_n51_n51# a_1237_1481#
X0 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X1 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X2 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X3 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X4 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X5 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X6 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X7 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X8 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X9 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X10 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X11 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X12 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X13 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X14 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X15 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X16 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X17 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X18 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X19 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X20 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X21 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X22 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X23 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X24 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X25 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X26 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X27 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X28 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X29 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X30 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X31 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X32 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X33 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X34 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X35 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X36 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X37 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X38 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X39 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X40 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X41 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X42 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X43 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X44 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
X45 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X46 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X47 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X48 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X49 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X50 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X51 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X52 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X53 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X54 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
X55 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
X56 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X57 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X58 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X59 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X60 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X61 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X62 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X63 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X64 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X65 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X66 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X67 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X68 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X69 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X70 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X71 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X72 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X73 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X74 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X75 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X76 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X77 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X78 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X79 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
.ends

.subckt comp018green_esd_rc_v5p0_1 VRC VPLUS VMINUS
X0 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X1 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X2 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X3 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X4 a_n2894_17198# a_n2614_4325# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X5 a_n1774_17198# a_n2054_4325# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X6 a_n1214_17198# a_n1494_4325# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X7 a_n2894_17198# a_n3174_4325# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X8 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X9 a_n2334_17198# a_n2614_4325# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X10 a_n1214_17198# a_n934_4325# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X11 a_n3454_17198# VPLUS VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X12 a_n1774_17198# a_n1494_4325# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X13 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X14 a_n2334_17198# a_n2054_4325# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X15 a_n654_17198# a_n934_4325# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X16 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X17 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X18 a_n3454_17198# a_n3174_4325# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X19 a_n654_17198# VRC VPLUS ppolyf_u r_width=0.8u r_length=63.855u
.ends

.subckt comp018green_esd_clamp_v5p0_1 top_route_0/VSUBS comp018green_esd_rc_v5p0_1_0/VPLUS
Xnmos_clamp_20_50_4_0 top_route_0/VSUBS comp018green_esd_rc_v5p0_1_0/VPLUS a_4685_27789#
+ nmos_clamp_20_50_4
Xcomp018green_esd_rc_v5p0_1_0 comp018green_esd_rc_v5p0_1_0/VRC comp018green_esd_rc_v5p0_1_0/VPLUS
+ top_route_0/VSUBS comp018green_esd_rc_v5p0_1
X0 a_2805_27789# comp018green_esd_rc_v5p0_1_0/VRC comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X1 comp018green_esd_rc_v5p0_1_0/VPLUS a_2805_27789# a_3781_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X2 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X3 a_3781_27789# a_2805_27789# top_route_0/VSUBS top_route_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X4 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X5 top_route_0/VSUBS a_3781_27789# a_4685_27789# top_route_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X6 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X7 comp018green_esd_rc_v5p0_1_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X8 a_4685_27789# a_3781_27789# top_route_0/VSUBS top_route_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X9 comp018green_esd_rc_v5p0_1_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X10 a_3781_27789# a_2805_27789# top_route_0/VSUBS top_route_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.7u
X11 top_route_0/VSUBS a_2805_27789# a_3781_27789# top_route_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X12 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.7u
X13 comp018green_esd_rc_v5p0_1_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X14 comp018green_esd_rc_v5p0_1_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X15 a_3781_27789# a_2805_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X16 comp018green_esd_rc_v5p0_1_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X17 top_route_0/VSUBS a_3781_27789# a_4685_27789# top_route_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X18 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X19 comp018green_esd_rc_v5p0_1_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X20 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X21 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X22 a_4685_27789# a_3781_27789# top_route_0/VSUBS top_route_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X23 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X24 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X25 a_2805_27789# comp018green_esd_rc_v5p0_1_0/VRC top_route_0/VSUBS top_route_0/VSUBS nfet_06v0 ad=2.2p pd=10.88u as=2.2p ps=10.88u w=5u l=0.7u
X26 comp018green_esd_rc_v5p0_1_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X27 top_route_0/VSUBS a_2805_27789# a_3781_27789# top_route_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X28 comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VRC a_2805_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X29 a_2805_27789# comp018green_esd_rc_v5p0_1_0/VRC comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.7u
X30 comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VRC a_2805_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X31 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X32 comp018green_esd_rc_v5p0_1_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X33 comp018green_esd_rc_v5p0_1_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X34 a_4685_27789# a_3781_27789# top_route_0/VSUBS top_route_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X35 top_route_0/VSUBS a_3781_27789# a_4685_27789# top_route_0/VSUBS nfet_06v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.7u
X36 comp018green_esd_rc_v5p0_1_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X37 comp018green_esd_rc_v5p0_1_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.7u
X38 a_3781_27789# a_2805_27789# top_route_0/VSUBS top_route_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X39 top_route_0/VSUBS a_2805_27789# a_3781_27789# top_route_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X40 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X41 a_3781_27789# a_2805_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.7u
X42 comp018green_esd_rc_v5p0_1_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X43 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_1_0/VPLUS comp018green_esd_rc_v5p0_1_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
.ends

.subckt comp018green_esd_clamp_v5p0_2 comp018green_esd_rc_v5p0_0/VPLUS top_route_1_0/VSUBS
Xnmos_clamp_20_50_4_0 top_route_1_0/VSUBS comp018green_esd_rc_v5p0_0/VPLUS a_4685_27789#
+ nmos_clamp_20_50_4
Xcomp018green_esd_rc_v5p0_0 comp018green_esd_rc_v5p0_0/VRC comp018green_esd_rc_v5p0_0/VPLUS
+ top_route_1_0/VSUBS comp018green_esd_rc_v5p0
X0 a_2805_27789# comp018green_esd_rc_v5p0_0/VRC comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X1 comp018green_esd_rc_v5p0_0/VPLUS a_2805_27789# a_3781_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X2 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X3 a_3781_27789# a_2805_27789# top_route_1_0/VSUBS top_route_1_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X4 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X5 top_route_1_0/VSUBS a_3781_27789# a_4685_27789# top_route_1_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X6 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X7 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X8 a_4685_27789# a_3781_27789# top_route_1_0/VSUBS top_route_1_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X9 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X10 a_3781_27789# a_2805_27789# top_route_1_0/VSUBS top_route_1_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.7u
X11 top_route_1_0/VSUBS a_2805_27789# a_3781_27789# top_route_1_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X12 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.7u
X13 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X14 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X15 a_3781_27789# a_2805_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X16 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X17 top_route_1_0/VSUBS a_3781_27789# a_4685_27789# top_route_1_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X18 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X19 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X20 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X21 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X22 a_4685_27789# a_3781_27789# top_route_1_0/VSUBS top_route_1_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X23 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X24 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X25 a_2805_27789# comp018green_esd_rc_v5p0_0/VRC top_route_1_0/VSUBS top_route_1_0/VSUBS nfet_06v0 ad=2.2p pd=10.88u as=2.2p ps=10.88u w=5u l=0.7u
X26 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X27 top_route_1_0/VSUBS a_2805_27789# a_3781_27789# top_route_1_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X28 comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VRC a_2805_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X29 a_2805_27789# comp018green_esd_rc_v5p0_0/VRC comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.7u
X30 comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VRC a_2805_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X31 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X32 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X33 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X34 a_4685_27789# a_3781_27789# top_route_1_0/VSUBS top_route_1_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X35 top_route_1_0/VSUBS a_3781_27789# a_4685_27789# top_route_1_0/VSUBS nfet_06v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.7u
X36 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X37 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.7u
X38 a_3781_27789# a_2805_27789# top_route_1_0/VSUBS top_route_1_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X39 top_route_1_0/VSUBS a_2805_27789# a_3781_27789# top_route_1_0/VSUBS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X40 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X41 a_3781_27789# a_2805_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.7u
X42 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27789# a_4685_27789# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X43 a_4685_27789# a_3781_27789# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
.ends

.subckt ESD_CLAMP_COR power_via_cor_3_0/m1_14757_49610# power_via_cor_5_0/m1_14757_35210#
+ power_via_cor_5_0/m1_14757_49610# comp018green_esd_clamp_v5p0_1_0/comp018green_esd_rc_v5p0_1_0/VPLUS
+ power_via_cor_3_0/m1_14757_35210# VSUBS comp018green_esd_clamp_v5p0_2_0/comp018green_esd_rc_v5p0_0/VPLUS
Xcomp018green_esd_clamp_v5p0_1_0 VSUBS comp018green_esd_clamp_v5p0_1_0/comp018green_esd_rc_v5p0_1_0/VPLUS
+ comp018green_esd_clamp_v5p0_1
Xcomp018green_esd_clamp_v5p0_2_0 comp018green_esd_clamp_v5p0_2_0/comp018green_esd_rc_v5p0_0/VPLUS
+ VSUBS comp018green_esd_clamp_v5p0_2
.ends

.subckt moscap_corner_2 VMINUS a_647_6541# a_5519_529#
X0 a_647_6541# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X1 a_5519_529# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X2 a_647_6541# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X3 a_5519_529# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X4 a_647_6541# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X5 a_647_6541# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
.ends

.subckt moscap_corner_3 VMINUS a_7955_529# a_3083_6541#
X0 a_7955_529# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X1 a_3083_6541# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X2 a_3083_6541# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X3 a_3083_6541# VMINUS cap_nmos_06v0 c_width=25u c_length=10u
.ends

.subckt GF_NI_COR_BASE VDD ESD_CLAMP_COR_0/power_via_cor_3_0/m1_14757_35210# ESD_CLAMP_COR_0/power_via_cor_3_0/m1_14757_49610#
+ ESD_CLAMP_COR_0/power_via_cor_5_0/m1_14757_35210# moscap_corner_0/a_647_6541# moscap_corner_6/a_647_529#
+ ESD_CLAMP_COR_0/power_via_cor_5_0/m1_14757_49610# moscap_corner_6/a_647_6541# moscap_corner_4/a_647_529#
+ moscap_corner_0/a_647_529# DVDD VSS moscap_corner_4/a_647_6541# moscap_corner_1/a_647_529#
Xmoscap_corner_1_0 moscap_corner_6/a_647_6541# moscap_corner_6/a_647_529# VSS moscap_corner_1
Xmoscap_corner_0 VSS moscap_corner_0/a_647_6541# moscap_corner_0/a_647_529# moscap_corner
Xmoscap_corner_1 VSS moscap_corner_1/a_647_529# moscap_corner_1/a_647_529# moscap_corner
Xmoscap_corner_2 VSS moscap_corner_4/a_647_6541# moscap_corner_4/a_647_529# moscap_corner
Xmoscap_corner_3 VSS moscap_corner_6/a_647_6541# moscap_corner_6/a_647_529# moscap_corner
Xmoscap_corner_5 VSS moscap_corner_6/a_647_6541# moscap_corner_6/a_647_529# moscap_corner
Xmoscap_corner_4 VSS moscap_corner_4/a_647_6541# moscap_corner_4/a_647_529# moscap_corner
Xmoscap_corner_6 VSS moscap_corner_6/a_647_6541# moscap_corner_6/a_647_529# moscap_corner
XESD_CLAMP_COR_0 ESD_CLAMP_COR_0/power_via_cor_3_0/m1_14757_49610# ESD_CLAMP_COR_0/power_via_cor_5_0/m1_14757_35210#
+ ESD_CLAMP_COR_0/power_via_cor_5_0/m1_14757_49610# VDD ESD_CLAMP_COR_0/power_via_cor_3_0/m1_14757_35210#
+ VSS DVDD ESD_CLAMP_COR
Xmoscap_corner_2_0 VSS moscap_corner_4/a_647_6541# moscap_corner_4/a_647_529# moscap_corner_2
Xmoscap_corner_3_0 VSS moscap_corner_1/a_647_529# moscap_corner_1/a_647_529# moscap_corner_3
.ends

.subckt gf180mcu_ocd_io__cor VDD DVDD VSS
XGF_NI_COR_BASE_0 VDD VSS VSS VSS DVDD DVDD VSS DVDD DVDD DVDD DVDD VSS DVDD DVDD
+ GF_NI_COR_BASE
.ends

.subckt GF_NI_VSS_BASE DVSS DVDD VDD m3_12861_12842# m3_7265_24036# m3_7265_54442#
+ m3_5168_44842# m3_9927_40042# m3_12297_28842# m3_7874_12842# m3_4851_11242# m3_7265_20836#
+ m3_7265_43242# m3_12297_24036# m3_12297_54442# m3_7265_41642# m3_4851_17636# m3_10244_48042#
+ m3_12297_20836# m3_2481_11242# m3_12297_43242# m3_12861_33636# m3_9927_28842# m3_12861_1636#
+ m3_12297_41642# m3_10244_44842# m3_2481_17636# m3_5168_1636# m3_12861_56043# m3_2798_27242#
+ m3_7874_33636# m3_9927_24036# m3_9927_54442# m3_7874_56043# m3_4851_30436# m3_7874_1636#
+ m3_9927_20836# m3_9927_43242# m3_2798_1636# m3_9927_41642# m3_7265_46442# m3_2798_12842#
+ m3_2481_30436# m3_7265_14436# m3_4851_40042# m3_5168_27242# m3_12861_8036# m3_5168_8036#
+ m3_12297_46442# m3_12861_4836# m3_12297_14436# m3_5168_4836# m3_2481_40042# m3_7874_8036#
+ m2_2292_38400# m3_12861_48042# m3_2798_8036# m3_4851_28842# m3_2798_33636# m3_5168_12842#
+ m3_7874_4836# m3_10244_1636# m3_9927_46442# m3_12861_44842# m3_7874_48042# m3_2798_56043#
+ m3_10244_27242# m3_4851_24036# m3_7265_11242# m3_2798_4836# m3_4851_54442# m3_9927_14436#
+ m3_2481_28842# m3_7874_44842# m3_7265_17636# m3_4851_20836# m3_4851_43242# m3_12297_11242#
+ m3_2481_24036# m3_2481_54442# m3_4851_41642# m3_5168_33636# m3_10244_12842# m3_12297_17636#
+ m3_2481_20836# m3_2481_43242# m3_10244_8036# m3_5168_56043# m3_2481_41642# m3_7265_30436#
+ m3_9927_11242# m3_10244_4836# m3_9927_17636# m3_2798_48042# m3_12297_30436# m3_10244_33636#
+ m3_7265_40042# m3_4851_46442# m3_2798_44842# m3_12861_27242# m3_10244_56043# m3_4851_14436#
+ VSS m3_12297_40042# m3_7874_27242# m3_2481_46442# comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS
+ m3_9927_30436# m3_2481_14436# m3_7265_28842# m3_5168_48042#
Xcomp018green_esd_clamp_v5p0_DVSS_0 comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS
+ VSS comp018green_esd_clamp_v5p0_DVSS
D0 VSS comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS diode_nd2ps_06v0 pj=82u area=40p
X0 comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS VSS cap_nmos_06v0 c_width=15u c_length=15u
D1 VSS comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS diode_nd2ps_06v0 pj=82u area=40p
D2 VSS comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS diode_nd2ps_06v0 pj=82u area=40p
D3 VSS comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS diode_nd2ps_06v0 pj=82u area=40p
X1 comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS VSS cap_nmos_06v0 c_width=15u c_length=15u
X2 comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS VSS cap_nmos_06v0 c_width=15u c_length=15u
X3 comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0/VPLUS VSS cap_nmos_06v0 c_width=15u c_length=15u
.ends

.subckt gf180mcu_ocd_io__vss VDD VSS DVDD DVSS
XGF_NI_VSS_BASE_0 DVSS DVDD VDD DVSS DVDD DVDD DVSS DVDD DVDD DVSS DVDD DVDD DVDD
+ DVDD DVDD DVDD DVDD DVSS DVDD DVDD DVDD DVSS DVDD DVSS DVDD DVSS DVDD DVSS DVSS
+ DVSS DVSS DVDD DVDD DVSS DVDD DVSS DVDD DVDD DVSS DVDD DVDD DVSS DVDD DVDD DVDD
+ DVSS DVSS DVSS DVDD DVSS DVDD DVSS DVDD DVSS VDD DVSS DVSS DVDD DVSS DVSS DVSS DVSS
+ DVDD DVSS DVSS DVSS DVSS DVDD DVDD DVSS DVDD DVDD DVDD DVSS DVDD DVDD DVDD DVDD
+ DVDD DVDD DVDD DVSS DVSS DVDD DVDD DVDD DVSS DVSS DVDD DVDD DVDD DVSS DVDD DVSS
+ DVDD DVSS DVDD DVDD DVSS DVSS DVSS DVDD VSS DVDD DVSS DVDD VDD DVDD DVDD DVDD DVSS
+ GF_NI_VSS_BASE
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_8 I ZN VDD VNW VPW VSS
X0 ZN I VDD VNW pfet_05v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1 VDD I ZN VNW pfet_05v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X2 ZN I VSS VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 ZN I VSS VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 ZN I VSS VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VDD I ZN VNW pfet_05v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X6 ZN I VDD VNW pfet_05v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X7 VSS I ZN VPW nfet_05v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 VDD I ZN VNW pfet_05v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X9 VSS I ZN VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X10 ZN I VDD VNW pfet_05v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X11 VSS I ZN VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X12 ZN I VDD VNW pfet_05v0 ad=0.4392p pd=1.94u as=0.5368p ps=3.32u w=1.22u l=0.5u
X13 VSS I ZN VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X14 ZN I VSS VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X15 VDD I ZN VNW pfet_05v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
D0 VPW I diode_nd2ps_06v0 pj=1.86u area=0.2052p
D1 I VNW diode_pd2nw_06v0 pj=1.86u area=0.2052p
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_12 I ZN VDD VNW VPW VSS
X0 ZN I VDD VNW pfet_05v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 ZN I VDD VNW pfet_05v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN I VSS VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 VSS I ZN VPW nfet_05v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 VDD I ZN VNW pfet_05v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5 ZN I VDD VNW pfet_05v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6 ZN I VSS VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7 ZN I VSS VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 VDD I ZN VNW pfet_05v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X9 ZN I VSS VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X10 ZN I VSS VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 VDD I ZN VNW pfet_05v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X12 VDD I ZN VNW pfet_05v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X13 ZN I VDD VNW pfet_05v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X14 VSS I ZN VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X15 VDD I ZN VNW pfet_05v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X16 VSS I ZN VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X17 VDD I ZN VNW pfet_05v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X18 VSS I ZN VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X19 ZN I VDD VNW pfet_05v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X20 VSS I ZN VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X21 ZN I VDD VNW pfet_05v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X22 VSS I ZN VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X23 ZN I VSS VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
X0 VDD a_572_375# a_484_472# VNW pfet_05v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VPW nfet_05v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VPW nfet_05v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 VDD a_124_375# a_36_472# VNW pfet_05v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
.ends

.subckt lvlshift_down VDD DVDD AH YL DVSS
Xgf180mcu_fd_sc_mcu7t5v0__inv_8_0 AH gf180mcu_fd_sc_mcu7t5v0__inv_8_0/ZN DVDD DVDD
+ DVSS DVSS gf180mcu_fd_sc_mcu7t5v0__inv_8
Xgf180mcu_fd_sc_mcu7t5v0__antenna_0 AH DVDD DVDD DVSS DVSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xgf180mcu_fd_sc_mcu7t5v0__inv_12_0 gf180mcu_fd_sc_mcu7t5v0__inv_8_0/ZN YL VDD VDD
+ DVSS DVSS gf180mcu_fd_sc_mcu7t5v0__inv_12
Xgf180mcu_fd_sc_mcu7t5v0__fillcap_8_0 DVDD DVDD DVSS DVSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
.ends

.subckt gf180mcu_ocd_io__fill10y VDD VSS AH YL DVDD DVSS
Xlvlshift_down_0 VDD DVDD AH YL DVSS lvlshift_down
XGF_NI_FILL10_0_0 DVSS DVDD VDD VSS GF_NI_FILL10_0short
.ends

.subckt GF_NI_FILL10_1pass VSS VDD DVSS DVDD m2_707_13108# m2_1290_13108#
XPOLY_SUB_FILL_1_0[0] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[1] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[2] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[3] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[4] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[5] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[6] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[7] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[8] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[9] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[10] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[11] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[12] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[13] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[14] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[15] VSS VDD POLY_SUB_FILL_1
.ends

.subckt GF_NI_FILL10_0pass DVSS DVDD VDD VSS GF_NI_FILL10_1_0/m2_1290_13108# GF_NI_FILL10_1_0/m2_707_13108#
XGF_NI_FILL10_1_0 VSS VDD DVSS DVDD GF_NI_FILL10_1_0/m2_707_13108# GF_NI_FILL10_1_0/m2_1290_13108#
+ GF_NI_FILL10_1pass
.ends

.subckt gf180mcu_ocd_io__fill10z DVDD DVSS VDD VSS thru0 thru1
XGF_NI_FILL10_0pass_0 DVSS DVDD VDD VSS thru1 thru0 GF_NI_FILL10_0pass
.ends

.subckt user_id_programming mask_rev[0] mask_rev[10] mask_rev[11] mask_rev[12] mask_rev[13]
+ mask_rev[14] mask_rev[15] mask_rev[16] mask_rev[17] mask_rev[18] mask_rev[19] mask_rev[1]
+ mask_rev[20] mask_rev[21] mask_rev[22] mask_rev[23] mask_rev[24] mask_rev[25] mask_rev[26]
+ mask_rev[27] mask_rev[28] mask_rev[29] mask_rev[2] mask_rev[30] mask_rev[31] mask_rev[3]
+ mask_rev[4] mask_rev[5] mask_rev[6] mask_rev[7] mask_rev[8] mask_rev[9] VDD VSS
Xmask_rev_value_one[9] VDD VDD VSS VSS mask_rev_value_one[9]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
XFILLCAP_4_3 VDD VDD VSS VSS gf180mcu_as_sc_mcu7t3v3__decap_4
Xmask_rev_value_one[8] VDD VDD VSS VSS mask_rev_value_one[8]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
XFILLCAP_4_4 VDD VDD VSS VSS gf180mcu_as_sc_mcu7t3v3__decap_4
Xmask_rev_value_one[7] VDD VDD VSS VSS mask_rev_value_one[7]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
XFILLCAP_4_5 VDD VDD VSS VSS gf180mcu_as_sc_mcu7t3v3__decap_4
Xmask_rev_value_one[6] VDD VDD VSS VSS mask_rev_value_one[6]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
XFILLCAP_4_6 VDD VDD VSS VSS gf180mcu_as_sc_mcu7t3v3__decap_4
Xmask_rev_value_one[5] VDD VDD VSS VSS mask_rev_value_one[5]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
XFILLCAP_4_7 VDD VDD VSS VSS gf180mcu_as_sc_mcu7t3v3__decap_4
Xmask_rev_value_one[4] VDD VDD VSS VSS mask_rev_value_one[4]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
XFILLCAP_4_8 VDD VDD VSS VSS gf180mcu_as_sc_mcu7t3v3__decap_4
Xmask_rev_value_one[3] VDD VDD VSS VSS mask_rev_value_one[3]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
XFILLCAP_4_9 VDD VDD VSS VSS gf180mcu_as_sc_mcu7t3v3__decap_4
Xmask_rev_value_one[19] VDD VDD VSS VSS mask_rev_value_one[19]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
Xmask_rev_value_one[2] VDD VDD VSS VSS mask_rev_value_one[2]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
Xmask_rev_value_one[18] VDD VDD VSS VSS mask_rev_value_one[18]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
Xmask_rev_value_one[1] VDD VDD VSS VSS mask_rev_value_one[1]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
Xmask_rev_value_one[17] VDD VDD VSS VSS mask_rev_value_one[17]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
Xmask_rev_value_one[0] VDD VDD VSS VSS mask_rev_value_one[0]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
Xmask_rev_value_one[16] VDD VDD VSS VSS mask_rev_value_one[16]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
Xmask_rev_value_zero[19] VDD VDD VSS VSS mask_rev[19] gf180mcu_as_sc_mcu7t3v3__tiel_4
Xmask_rev_value_one[15] VDD VDD VSS VSS mask_rev_value_one[15]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
Xmask_rev_value_one[31] VDD VDD VSS VSS mask_rev_value_one[31]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
Xmask_rev_value_zero[18] VDD VDD VSS VSS mask_rev[18] gf180mcu_as_sc_mcu7t3v3__tiel_4
Xmask_rev_value_one[14] VDD VDD VSS VSS mask_rev_value_one[14]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
Xmask_rev_value_one[30] VDD VDD VSS VSS mask_rev_value_one[30]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
Xmask_rev_value_zero[17] VDD VDD VSS VSS mask_rev[17] gf180mcu_as_sc_mcu7t3v3__tiel_4
Xmask_rev_value_one[13] VDD VDD VSS VSS mask_rev_value_one[13]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
Xmask_rev_value_zero[16] VDD VDD VSS VSS mask_rev[16] gf180mcu_as_sc_mcu7t3v3__tiel_4
Xmask_rev_value_one[12] VDD VDD VSS VSS mask_rev_value_one[12]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
Xmask_rev_value_zero[15] VDD VDD VSS VSS mask_rev[15] gf180mcu_as_sc_mcu7t3v3__tiel_4
Xmask_rev_value_one[11] VDD VDD VSS VSS mask_rev_value_one[11]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
XFILLCAP_4_20 VDD VDD VSS VSS gf180mcu_as_sc_mcu7t3v3__decap_4
Xmask_rev_value_zero[31] VDD VDD VSS VSS mask_rev[31] gf180mcu_as_sc_mcu7t3v3__tiel_4
Xmask_rev_value_one[10] VDD VDD VSS VSS mask_rev_value_one[10]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
Xmask_rev_value_zero[14] VDD VDD VSS VSS mask_rev[14] gf180mcu_as_sc_mcu7t3v3__tiel_4
XFILLCAP_4_21 VDD VDD VSS VSS gf180mcu_as_sc_mcu7t3v3__decap_4
Xmask_rev_value_zero[30] VDD VDD VSS VSS mask_rev[30] gf180mcu_as_sc_mcu7t3v3__tiel_4
XFILLCAP_4_10 VDD VDD VSS VSS gf180mcu_as_sc_mcu7t3v3__decap_4
Xmask_rev_value_zero[13] VDD VDD VSS VSS mask_rev[13] gf180mcu_as_sc_mcu7t3v3__tiel_4
XFILLCAP_4_22 VDD VDD VSS VSS gf180mcu_as_sc_mcu7t3v3__decap_4
XFILLCAP_4_11 VDD VDD VSS VSS gf180mcu_as_sc_mcu7t3v3__decap_4
Xmask_rev_value_zero[12] VDD VDD VSS VSS mask_rev[12] gf180mcu_as_sc_mcu7t3v3__tiel_4
XFILLCAP_4_23 VDD VDD VSS VSS gf180mcu_as_sc_mcu7t3v3__decap_4
XFILLCAP_4_12 VDD VDD VSS VSS gf180mcu_as_sc_mcu7t3v3__decap_4
Xmask_rev_value_zero[11] VDD VDD VSS VSS mask_rev[11] gf180mcu_as_sc_mcu7t3v3__tiel_4
Xmask_rev_value_zero[9] VDD VDD VSS VSS mask_rev[9] gf180mcu_as_sc_mcu7t3v3__tiel_4
XFILLCAP_4_13 VDD VDD VSS VSS gf180mcu_as_sc_mcu7t3v3__decap_4
Xmask_rev_value_zero[8] VDD VDD VSS VSS mask_rev[8] gf180mcu_as_sc_mcu7t3v3__tiel_4
Xmask_rev_value_zero[10] VDD VDD VSS VSS mask_rev[10] gf180mcu_as_sc_mcu7t3v3__tiel_4
XFILLCAP_4_14 VDD VDD VSS VSS gf180mcu_as_sc_mcu7t3v3__decap_4
Xmask_rev_value_zero[7] VDD VDD VSS VSS mask_rev[7] gf180mcu_as_sc_mcu7t3v3__tiel_4
XFILLCAP_4_15 VDD VDD VSS VSS gf180mcu_as_sc_mcu7t3v3__decap_4
Xmask_rev_value_zero[6] VDD VDD VSS VSS mask_rev[6] gf180mcu_as_sc_mcu7t3v3__tiel_4
XFILLCAP_4_16 VDD VDD VSS VSS gf180mcu_as_sc_mcu7t3v3__decap_4
Xmask_rev_value_zero[5] VDD VDD VSS VSS mask_rev[5] gf180mcu_as_sc_mcu7t3v3__tiel_4
XFILLCAP_4_17 VDD VDD VSS VSS gf180mcu_as_sc_mcu7t3v3__decap_4
Xmask_rev_value_one[29] VDD VDD VSS VSS mask_rev_value_one[29]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
Xmask_rev_value_zero[4] VDD VDD VSS VSS mask_rev[4] gf180mcu_as_sc_mcu7t3v3__tiel_4
XFILLCAP_4_18 VDD VDD VSS VSS gf180mcu_as_sc_mcu7t3v3__decap_4
Xmask_rev_value_one[28] VDD VDD VSS VSS mask_rev_value_one[28]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
Xmask_rev_value_zero[3] VDD VDD VSS VSS mask_rev[3] gf180mcu_as_sc_mcu7t3v3__tiel_4
XFILLCAP_4_19 VDD VDD VSS VSS gf180mcu_as_sc_mcu7t3v3__decap_4
Xmask_rev_value_one[27] VDD VDD VSS VSS mask_rev_value_one[27]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
Xmask_rev_value_zero[2] VDD VDD VSS VSS mask_rev[2] gf180mcu_as_sc_mcu7t3v3__tiel_4
Xmask_rev_value_one[26] VDD VDD VSS VSS mask_rev_value_one[26]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
Xmask_rev_value_zero[1] VDD VDD VSS VSS mask_rev[1] gf180mcu_as_sc_mcu7t3v3__tiel_4
Xmask_rev_value_zero[29] VDD VDD VSS VSS mask_rev[29] gf180mcu_as_sc_mcu7t3v3__tiel_4
Xmask_rev_value_one[25] VDD VDD VSS VSS mask_rev_value_one[25]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
Xmask_rev_value_zero[0] VDD VDD VSS VSS mask_rev[0] gf180mcu_as_sc_mcu7t3v3__tiel_4
Xmask_rev_value_zero[28] VDD VDD VSS VSS mask_rev[28] gf180mcu_as_sc_mcu7t3v3__tiel_4
Xmask_rev_value_one[24] VDD VDD VSS VSS mask_rev_value_one[24]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
Xmask_rev_value_zero[27] VDD VDD VSS VSS mask_rev[27] gf180mcu_as_sc_mcu7t3v3__tiel_4
Xmask_rev_value_one[23] VDD VDD VSS VSS mask_rev_value_one[23]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
Xmask_rev_value_zero[26] VDD VDD VSS VSS mask_rev[26] gf180mcu_as_sc_mcu7t3v3__tiel_4
Xmask_rev_value_one[22] VDD VDD VSS VSS mask_rev_value_one[22]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
Xmask_rev_value_zero[25] VDD VDD VSS VSS mask_rev[25] gf180mcu_as_sc_mcu7t3v3__tiel_4
Xmask_rev_value_one[21] VDD VDD VSS VSS mask_rev_value_one[21]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
Xmask_rev_value_zero[24] VDD VDD VSS VSS mask_rev[24] gf180mcu_as_sc_mcu7t3v3__tiel_4
Xmask_rev_value_one[20] VDD VDD VSS VSS mask_rev_value_one[20]/ONE gf180mcu_as_sc_mcu7t3v3__tieh_4
Xmask_rev_value_zero[23] VDD VDD VSS VSS mask_rev[23] gf180mcu_as_sc_mcu7t3v3__tiel_4
XFILLCAP_4_0 VDD VDD VSS VSS gf180mcu_as_sc_mcu7t3v3__decap_4
Xmask_rev_value_zero[22] VDD VDD VSS VSS mask_rev[22] gf180mcu_as_sc_mcu7t3v3__tiel_4
XFILLCAP_4_1 VDD VDD VSS VSS gf180mcu_as_sc_mcu7t3v3__decap_4
Xmask_rev_value_zero[21] VDD VDD VSS VSS mask_rev[21] gf180mcu_as_sc_mcu7t3v3__tiel_4
XFILLCAP_4_2 VDD VDD VSS VSS gf180mcu_as_sc_mcu7t3v3__decap_4
Xmask_rev_value_zero[20] VDD VDD VSS VSS mask_rev[20] gf180mcu_as_sc_mcu7t3v3__tiel_4
.ends

.subckt tie_poly_res a_n2051_55943# a_n2051_55061# a_n2331_55943# w_n2756_54700#
X0 a_n2051_55943# a_n2051_55061# w_n2756_54700# ppolyf_u r_width=0.8u r_length=3.9u
X1 a_n2331_55943# w_n2756_54700# w_n2756_54700# ppolyf_u r_width=0.8u r_length=3.9u
.ends

.subckt GF_NI_IN_S_BASE PD PU Y ndrive_y_<0> ndrive_x_<0> ndrive_x_<1> ndrive_Y_<1>
+ ndrive_x_<2> ndrive_y_<2> ndrive_x_<3> ndrive_Y_<3> pdrive_x_<0> pdrive_y_<0> pdrive_y_<1>
+ pdrive_x_<1> pdrive_x_<2> pdrive_y_<2> pdrive_y_<3> pdrive_x_<3> m3_1771_39126#
+ w_11000_43887# comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_4/m1_n44_0#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/w_n5_111#
+ m2_1886_52816# comp018green_inpath_cms_smt_0/m3_9619_4882# w_835_53274# comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_1/m1_n44_400#
+ comp018green_inpath_cms_smt_0/m3_9619_3696# comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_2/m1_n44_400#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_3/m1_n44_400#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_5/m1_n44_0#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_1/m1_n44_0#
+ comp018green_esd_cdm_0/w_454_3720# m3_10025_37504# PAD comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_2/m1_n44_0#
+ a_12390_41548# m1_3608_46684# comp018green_esd_cdm_0/DVDD comp018green_inpath_cms_smt_0/comp018green_sigbuf_3/DVDD
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_3/m1_n44_0#
+ tie_poly_res_0/VSUBS comp018green_sigbuf_1_0/DVSS comp018green_esd_cdm_0/DVSS comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VDD
+ comp018green_sigbuf_1_0/DVDD comp018green_inpath_cms_smt_0/m1_10570_5335# comp018green_inpath_cms_smt_0/VSUBS
+ w_11042_41027# comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/VSUBS
+ comp018green_out_predrv_3/DVDD w_13720_39292# comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS
Xlv_nand_2 tie_poly_res_0/VSUBS w_13720_39292# w_11184_44921# m1_5236_36986# w_13720_39292#
+ lv_nand
Xlv_nand_3 tie_poly_res_0/VSUBS w_13720_39292# w_11184_44921# m1_4812_38523# w_11184_44921#
+ lv_nand
Xcomp018green_out_paddrv_16T_0 pdrive_x_<2> pdrive_x_<3> pdrive_y_<3> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_4/m1_n44_0#
+ pdrive_x_<3> ndrive_Y_<3> pdrive_x_<0> pdrive_x_<2> pdrive_y_<0> comp018green_out_predrv_3/DVDD
+ ndrive_x_<0> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/w_n5_111#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_1/m1_n44_0#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_5/m1_n44_0#
+ ndrive_y_<2> pdrive_y_<2> pdrive_x_<1> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_1/m1_n44_400#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_2/m1_n44_400#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_3/m1_n44_400#
+ ndrive_x_<3> pdrive_y_<1> ndrive_x_<1> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_2/m1_n44_0#
+ ndrive_y_<0> pdrive_x_<0> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/VSUBS
+ ndrive_x_<2> pdrive_x_<1> PAD ndrive_Y_<1> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_3/m1_n44_0#
+ comp018green_out_paddrv_16T
Xtie_poly_res_0 w_11184_44921# comp018green_inpath_cms_smt_0/VSUBS comp018green_inpath_cms_smt_0/CS
+ w_835_53274# tie_poly_res
Xcomp018green_sigbuf_1_0 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/DVSS comp018green_sigbuf_1_0/DVDD
+ comp018green_sigbuf_1_0/ZB m1_9774_36986# m1_9537_37107# comp018green_sigbuf_1
Xcomp018green_out_predrv_0 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/ZB ndrive_x_<0>
+ comp018green_out_predrv_0/ENB comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_3/A
+ comp018green_out_predrv_3/DVDD ndrive_y_<0> pdrive_y_<0> pdrive_x_<0> comp018green_out_predrv_0/EN
+ comp018green_out_predrv
Xcomp018green_out_sigbuf_a_0 comp018green_out_predrv_3/A comp018green_sigbuf_1_0/DVSS
+ comp018green_sigbuf_1_0/DVDD m1_9174_38525# m1_9257_38818# comp018green_out_sigbuf_a
Xcomp018green_out_predrv_2 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/ZB ndrive_x_<2>
+ comp018green_out_predrv_3/ENB comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_3/A
+ comp018green_out_predrv_3/DVDD ndrive_y_<2> pdrive_y_<2> pdrive_x_<2> comp018green_out_predrv_3/EN
+ comp018green_out_predrv
Xcomp018green_out_predrv_1 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/ZB ndrive_x_<3>
+ comp018green_out_predrv_1/ENB comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_3/A
+ comp018green_out_predrv_3/DVDD ndrive_Y_<3> pdrive_y_<3> pdrive_x_<3> comp018green_out_predrv_1/EN
+ comp018green_out_predrv
Xcomp018green_out_sigbuf_oe_0 comp018green_out_predrv_0/ENB comp018green_sigbuf_1_0/DVDD
+ comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_0/EN m1_1178_38534# m1_1183_38806#
+ comp018green_out_sigbuf_oe
Xcomp018green_out_predrv_3 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/ZB ndrive_x_<1>
+ comp018green_out_predrv_3/ENB comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_3/A
+ comp018green_out_predrv_3/DVDD ndrive_Y_<1> pdrive_y_<1> pdrive_x_<1> comp018green_out_predrv_3/EN
+ comp018green_out_predrv
Xcomp018green_inpath_cms_smt_0 comp018green_esd_cdm_0/IP_IN comp018green_inpath_cms_smt_0/CS
+ PU comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VDD comp018green_inpath_cms_smt_0/CS
+ w_11000_43887# m1_3608_46684# comp018green_esd_cdm_0/IP_IN comp018green_inpath_cms_smt_0/m3_9619_4882#
+ comp018green_inpath_cms_smt_0/m3_9619_3696# comp018green_esd_cdm_0/DVSS comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VDD
+ comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS
+ Y comp018green_inpath_cms_smt_0/VSUBS comp018green_inpath_cms_smt_0/m1_10570_5335#
+ comp018green_inpath_cms_smt_0/comp018green_in_pupd_0/a_506_484# PD w_835_53274#
+ comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS comp018green_inpath_cms_smt_0/comp018green_sigbuf_3/DVDD
+ comp018green_inpath_cms_smt
Xcomp018green_out_sigbuf_oe_2 comp018green_out_predrv_1/ENB comp018green_sigbuf_1_0/DVDD
+ comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_1/EN m1_5236_36986# m1_5084_37107#
+ comp018green_out_sigbuf_oe
Xcomp018green_out_sigbuf_oe_1 comp018green_out_predrv_3/ENB comp018green_sigbuf_1_0/DVDD
+ comp018green_sigbuf_1_0/DVSS comp018green_out_predrv_3/EN m1_4812_38523# m1_4626_36747#
+ comp018green_out_sigbuf_oe
Xlv_inv_0 w_13720_39292# m1_1183_38806# m1_1178_38534# tie_poly_res_0/VSUBS lv_inv
Xlv_inv_1 w_13720_39292# m1_9257_38818# m1_9174_38525# tie_poly_res_0/VSUBS lv_inv
Xlv_inv_2 w_13720_39292# m1_9537_37107# m1_9774_36986# tie_poly_res_0/VSUBS lv_inv
Xlv_inv_3 w_13720_39292# m1_4626_36747# m1_4812_38523# tie_poly_res_0/VSUBS lv_inv
Xlv_inv_4 w_13720_39292# m1_9774_36986# w_11184_44921# tie_poly_res_0/VSUBS lv_inv
Xlv_inv_6 w_13720_39292# m1_5084_37107# m1_5236_36986# tie_poly_res_0/VSUBS lv_inv
Xcomp018green_esd_cdm_0 comp018green_esd_cdm_0/IP_IN PAD comp018green_esd_cdm_0/DVDD
+ comp018green_esd_cdm_0/DVSS comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VDD
+ comp018green_esd_cdm_0/w_454_3720# comp018green_esd_cdm
Xlv_nand_0 tie_poly_res_0/VSUBS w_13720_39292# w_11184_44921# m1_9174_38525# w_11184_44921#
+ lv_nand
Xlv_nand_1 tie_poly_res_0/VSUBS w_13720_39292# w_11184_44921# m1_1178_38534# w_11184_44921#
+ lv_nand
X0 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X1 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X2 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X3 a_12390_41548# comp018green_esd_cdm_0/DVSS cap_nmos_06v0 c_width=3u c_length=3u
X4 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X5 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X6 a_12390_41548# comp018green_esd_cdm_0/DVSS cap_nmos_06v0 c_width=3u c_length=3u
X7 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
X8 a_12390_41548# comp018green_esd_cdm_0/DVSS cap_nmos_06v0 c_width=3u c_length=3u
X9 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
D0 comp018green_inpath_cms_smt_0/VSUBS w_11184_44921# diode_pd2nw_03v3 pj=1.92u area=0.2304p
D1 comp018green_inpath_cms_smt_0/VSUBS w_11184_44921# diode_pd2nw_03v3 pj=1.92u area=0.2304p
D2 comp018green_inpath_cms_smt_0/VSUBS w_11184_44921# diode_pd2nw_03v3 pj=1.92u area=0.2304p
D3 comp018green_inpath_cms_smt_0/VSUBS w_11000_43887# diode_pd2nw_03v3 pj=1.92u area=0.2304p
D4 w_11184_44921# w_11042_41027# diode_pd2nw_03v3 pj=4u area=1p
D5 w_11184_44921# w_11042_41027# diode_pd2nw_03v3 pj=4u area=1p
X10 a_12390_41548# comp018green_esd_cdm_0/DVSS cap_nmos_06v0 c_width=3u c_length=3u
D6 comp018green_inpath_cms_smt_0/VSUBS w_11184_44921# diode_pd2nw_03v3 pj=1.92u area=0.2304p
D7 comp018green_inpath_cms_smt_0/VSUBS w_11184_44921# diode_pd2nw_03v3 pj=1.92u area=0.2304p
X11 comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/VSS cap_nmos_06v0 c_width=5u c_length=1.5u
.ends

.subckt gf180mcu_ocd_io__in_s DVDD PD PU VDD PAD Y VSS DVSS
XGF_NI_IN_S_BASE_0 PD PU Y GF_NI_IN_S_BASE_0/ndrive_y_<0> GF_NI_IN_S_BASE_0/ndrive_x_<0>
+ GF_NI_IN_S_BASE_0/ndrive_x_<1> GF_NI_IN_S_BASE_0/ndrive_Y_<1> GF_NI_IN_S_BASE_0/ndrive_x_<2>
+ GF_NI_IN_S_BASE_0/ndrive_y_<2> GF_NI_IN_S_BASE_0/ndrive_x_<3> GF_NI_IN_S_BASE_0/ndrive_Y_<3>
+ GF_NI_IN_S_BASE_0/pdrive_x_<0> GF_NI_IN_S_BASE_0/pdrive_y_<0> GF_NI_IN_S_BASE_0/pdrive_y_<1>
+ GF_NI_IN_S_BASE_0/pdrive_x_<1> GF_NI_IN_S_BASE_0/pdrive_x_<2> GF_NI_IN_S_BASE_0/pdrive_y_<2>
+ GF_NI_IN_S_BASE_0/pdrive_y_<3> GF_NI_IN_S_BASE_0/pdrive_x_<3> VDD VDD DVDD DVDD
+ DVSS VDD VDD DVSS VSS DVSS DVSS DVDD DVDD DVDD VSS PAD DVDD DVDD DVDD DVDD DVDD
+ DVDD VSS DVSS DVSS DVDD DVDD VDD VSS VDD DVSS DVDD VDD DVSS GF_NI_IN_S_BASE
.ends

.subckt gf180mcu_padframe gpio_in[38] gpio[39] gpio_in[39] gpio_drive2[38] gpio_in[43]
+ gpio[10] gpio[13] gpio[16] gpio[19] gpio[22] gpio[25] gpio[2] gpio[30] gpio[32]
+ gpio[33] gpio[35] gpio[36] gpio_drive0[0] gpio_drive0[5] gpio_drive1[6] gpio_drive1[7]
+ gpio_drive1[8] gpio_drive0[9] gpio_drive1[9] gpio_drive0[10] gpio_drive0[11] gpio_drive0[12]
+ gpio_drive0[13] gpio_drive1[13] gpio_drive0[14] gpio_drive0[1] gpio_drive0[15] gpio_drive0[16]
+ gpio_drive0[17] gpio_drive0[18] gpio_drive1[18] gpio_drive1[1] gpio_drive1[21] gpio_drive1[22]
+ gpio_drive0[23] gpio_drive1[23] gpio_drive0[24] gpio_drive1[24] gpio_drive0[2] gpio_drive1[26]
+ gpio_drive1[27] gpio_drive0[28] gpio_drive1[28] gpio_drive0[29] gpio_drive1[29]
+ gpio_drive1[2] gpio_drive1[30] gpio_drive0[32] gpio_drive0[33] gpio_drive0[34] gpio_drive0[3]
+ gpio_drive0[35] gpio_drive1[35] gpio_drive0[36] gpio_drive1[3] gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[29]
+ gpio_in[2] gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[34] gpio_in[35]
+ gpio_in[36] gpio_in[37] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_ie[10] gpio_ie[11] gpio_ie[12] gpio_ie[13] gpio_ie[14] gpio_ie[24] gpio_ie[25]
+ gpio_ie[28] gpio_ie[29] gpio_ie[2] gpio_ie[30] gpio_ie[33] gpio_ie[5] gpio_ie[6]
+ gpio_ie[9] gpio_out[10] gpio_out[11] gpio_out[13] gpio_out[14] gpio_out[17] gpio_out[19]
+ gpio_out[22] gpio_out[25] gpio_out[28] gpio_out[30] gpio_out[32] gpio_out[33] gpio_out[34]
+ gpio_out[35] gpio_out[36] gpio_out[37] gpio_out[6] gpio_out[9] gpio_oe[10] gpio_oe[12]
+ gpio_oe[13] gpio_oe[15] gpio_oe[16] gpio_oe[17] gpio_oe[18] gpio_oe[19] gpio_oe[24]
+ gpio_oe[27] gpio_oe[28] gpio_oe[30] gpio_oe[31] gpio_oe[33] gpio_oe[34] gpio_oe[35]
+ gpio_oe[36] gpio_oe[8] gpio_pulldown[11] gpio_pulldown[15] gpio_pulldown[1] gpio_pulldown[21]
+ gpio_pulldown[22] gpio_pulldown[24] gpio_pulldown[25] gpio_pulldown[27] gpio_pulldown[28]
+ gpio_pulldown[29] gpio_pulldown[2] gpio_pulldown[33] gpio_pulldown[36] gpio_pulldown[5]
+ gpio_pulldown[8] gpio_pulldown[9] gpio_pullup[0] gpio_pullup[10] gpio_pullup[11]
+ gpio_pullup[12] gpio_pullup[13] gpio_pullup[14] gpio_pullup[15] gpio_pullup[1] gpio_pullup[25]
+ gpio_pullup[26] gpio_pullup[28] gpio_pullup[29] gpio_pullup[30] gpio_pullup[31]
+ gpio_pullup[32] gpio_pullup[33] gpio_pullup[37] gpio_pullup[3] gpio_pullup[4] gpio_pullup[6]
+ gpio_pullup[7] gpio_pullup[8] gpio_pullup[9] gpio_schmitt[11] gpio_schmitt[12] gpio_schmitt[13]
+ gpio_schmitt[14] gpio_schmitt[15] gpio_schmitt[1] gpio_schmitt[20] gpio_schmitt[24]
+ gpio_schmitt[26] gpio_schmitt[27] gpio_schmitt[29] gpio_schmitt[2] gpio_schmitt[30]
+ gpio_schmitt[31] gpio_schmitt[32] gpio_schmitt[4] gpio_schmitt[5] gpio_schmitt[6]
+ gpio_schmitt[7] gpio_schmitt[8] gpio_schmitt[9] gpio_slew[0] gpio_slew[15] gpio_slew[22]
+ gpio_slew[24] gpio_slew[25] gpio_slew[26] gpio_slew[27] gpio_slew[28] gpio_slew[29]
+ gpio_slew[2] gpio_slew[33] gpio_slew[36] gpio_slew[3] gpio_slew[4] gpio_slew[5]
+ gpio_slew[6] gpio_slew[7] gpio_slew[8] gpio_slew[9] resetb_core gpio_ana[0] gpio_ana[1]
+ gpio_ana[2] gpio_ana[3] gpio_ana[4] gpio_ana[5] gpio_ana[6] gpio_ana[7] gpio_ana[8]
+ gpio_ana[9] gpio_ana[10] gpio_ana[11] gpio_ana[12] gpio_ana[13] gpio_ana[14] gpio_ana[18]
+ gpio_ana[21] gpio_ana[22] gpio_ana[23] gpio_ana[24] gpio_ana[25] gpio_ana[26] gpio_ana[27]
+ gpio_ana[28] gpio_ana[29] gpio_ana[30] gpio_ana[31] gpio_ana[32] gpio_ana[33] gpio_ana[34]
+ gpio_ana[35] gpio_ana[36] gpio_ana[37] gpio_ana[40] gpio_ana[41] gpio_ana[42] gpio_ana[43]
+ gpio_loopback_zero[0] gpio_loopback_one[0] gpio_loopback_zero[1] gpio_loopback_one[1]
+ gpio_loopback_zero[2] gpio_loopback_one[2] gpio_loopback_one[3] gpio_loopback_zero[3]
+ gpio_loopback_zero[4] gpio_loopback_one[4] gpio_loopback_one[5] gpio_loopback_zero[5]
+ gpio_loopback_zero[6] gpio_loopback_one[6] gpio_loopback_one[7] gpio_loopback_zero[7]
+ gpio_loopback_zero[8] gpio_loopback_one[8] gpio_loopback_one[9] gpio_loopback_zero[9]
+ gpio_loopback_zero[10] gpio_loopback_one[11] gpio_loopback_zero[11] gpio_loopback_zero[12]
+ gpio_loopback_one[12] gpio_loopback_one[13] gpio_loopback_zero[14] gpio_loopback_one[14]
+ gpio_loopback_one[15] gpio_loopback_zero[15] gpio_loopback_zero[16] gpio_loopback_one[16]
+ gpio_loopback_one[17] gpio_loopback_zero[17] gpio_loopback_zero[18] gpio_loopback_one[18]
+ gpio_loopback_one[19] gpio_loopback_zero[19] gpio_loopback_zero[20] gpio_loopback_one[20]
+ gpio_loopback_one[21] gpio_loopback_zero[21] gpio_loopback_one[22] gpio_loopback_one[23]
+ gpio_loopback_zero[23] gpio_loopback_zero[24] gpio_loopback_one[25] gpio_loopback_zero[25]
+ gpio_loopback_zero[26] gpio_loopback_one[26] gpio_loopback_one[27] gpio_loopback_zero[27]
+ gpio_loopback_zero[28] gpio_loopback_one[28] gpio_loopback_one[29] gpio_loopback_zero[29]
+ gpio_loopback_zero[30] gpio_loopback_one[30] gpio_loopback_one[31] gpio_loopback_zero[31]
+ gpio_loopback_zero[32] gpio_loopback_one[32] gpio_loopback_zero[33] gpio_loopback_zero[34]
+ gpio_loopback_one[34] gpio_loopback_one[35] gpio_loopback_zero[35] gpio_loopback_zero[36]
+ gpio_loopback_one[36] gpio_loopback_one[37] gpio_loopback_zero[37] gpio_loopback_zero[38]
+ gpio_loopback_zero[39] gpio_loopback_zero[40] gpio_loopback_one[40] gpio_loopback_one[41]
+ gpio_loopback_one[43] gpio_loopback_zero[43] resetb_loopback_zero porb_h porb_l
+ mask_rev[0] mask_rev[1] mask_rev[2] mask_rev[3] mask_rev[4] mask_rev[5] mask_rev[6]
+ mask_rev[7] mask_rev[8] mask_rev[9] mask_rev[20] mask_rev[21] mask_rev[22] mask_rev[23]
+ mask_rev[24] mask_rev[25] mask_rev[26] gpio_drive0[30] gpio_drive0[42] gpio_drive1[42]
+ gpio_pulldown[42] gpio_pullup[41] gpio_drive0[41] gpio_drive1[41] gpio_slew[41]
+ gpio_schmitt[40] gpio_out[39] gpio_oe[43] gpio_slew[43] gpio_ie[43] gpio_pulldown[43]
+ gpio_drive1[43] gpio_ie[15] gpio_pullup[34] gpio_schmitt[35] gpio_out[3] gpio_out[0]
+ gpio_loopback_one[10] gpio_drive1[12] gpio_oe[5] gpio_slew[12] gpio_slew[30] gpio_ie[37]
+ gpio_ana[15] gpio_oe[2] gpio_drive0[8] gpio_drive1[17] gpio_pullup[38] resetb_loopback_one
+ gpio_pulldown[12] gpio_drive1[34] gpio_pulldown[30] gpio_ie[16] gpio_ie[34] gpio_loopback_one[33]
+ gpio_slew[37] gpio_drive1[11] mask_rev[27] gpio[0] gpio_pullup[17] mask_rev[29]
+ gpio_in[20] gpio_schmitt[18] gpio_pullup[35] gpio_schmitt[36] gpio[23] gpio_out[8]
+ gpio_ie[3] gpio_oe[9] gpio_slew[16] gpio_ie[31] mask_rev[28] gpio_slew[34] gpio_out[5]
+ gpio[3] gpio_oe[37] gpio_slew[39] mask_rev[31] gpio_out[27] gpio_drive0[38] gpio_out[2]
+ gpio_out[24] gpio_in[40] gpio_drive0[7] gpio_in[28] mask_rev[30] gpio_drive0[22]
+ gpio_in[22] gpio_drive1[16] gpio[42] gpio_oe[42] gpio_schmitt[33] gpio_pulldown[19]
+ gpio[20] gpio_pulldown[37] gpio_ie[0] por_h gpio_oe[6] gpio_slew[13] gpio_ana[19]
+ gpio_slew[31] gpio_oe[25] gpio_oe[39] gpio_drive1[33] gpio[41] gpio_loopback_zero[22]
+ mask_rev[11] gpio_drive1[10] gpio_ie[38] gpio[43] gpio_drive0[43] gpio[26] gpio_pulldown[6]
+ gpio_pullup[20] gpio_pullup[19] gpio_pullup[40] gpio_schmitt[21] gpio_pulldown[16]
+ gpio_out[21] gpio_pulldown[34] gpio_ie[41] mask_rev[10] gpio_pulldown[39] gpio_drive0[27]
+ mask_rev[13] gpio_ana[16] gpio_oe[3] gpio[6] gpio_slew[10] gpio_oe[22] gpio_schmitt[43]
+ mask_rev[12] gpio_pullup[42] gpio_loopback_one[38] mask_rev[15] gpio_schmitt[23]
+ gpio_slew[38] gpio_drive0[6] gpio_pulldown[3] gpio_pulldown[13] mask_rev[14] gpio_ie[7]
+ gpio_drive0[21] gpio_pulldown[31] gpio_ie[17] gpio_drive1[15] gpio_ie[26] mask_rev[17]
+ gpio_ie[35] gpio_drive1[39] gpio_out[41] gpio_oe[0] gpio_drive1[0] mask_rev[16]
+ gpio_drive0[39] gpio_in[6] mask_rev[19] gpio[1] gpio_out[42] gpio_drive1[32] gpio_slew[18]
+ gpio_loopback_zero[41] gpio_pullup[18] gpio_pullup[27] gpio_schmitt[19] gpio_pullup[36]
+ gpio_schmitt[28] gpio_schmitt[37] gpio[29] mask_rev[18] gpio_oe[38] gpio_pulldown[0]
+ gpio_pulldown[10] gpio_ie[4] resetb_pullup gpio_ie[23] gpio_pullup[22] gpio_ie[32]
+ gpio_slew[17] gpio_oe[41] gpio_slew[35] gpio_oe[29] gpio[9] gpio_pullup[39] gpio[14]
+ gpio_out[43] gpio_out[7] gpio_drive0[26] gpio_out[29] gpio[11] resetb_pulldown gpio_schmitt[42]
+ gpio_ana[20] gpio_out[4] gpio_pulldown[38] gpio_out[26] gpio_loopback_zero[42] gpio_pullup[5]
+ gpio_out[31] gpio_drive1[5] gpio_pullup[24] gpio_ie[21] gpio_schmitt[16] gpio_out[1]
+ gpio_pulldown[41] gpio[24] gpio_schmitt[25] gpio[40] gpio_schmitt[34] gpio[21] gpio_out[23]
+ gpio_loopback_one[24] gpio_loopback_zero[13] gpio_schmitt[39] gpio_drive1[20] gpio_ie[1]
+ gpio_drive1[37] gpio_out[15] gpio_ie[20] gpio_ie[19] gpio_oe[7] gpio_slew[14] gpio_ie[40]
+ gpio_slew[23] gpio_out[20] gpio[4] gpio_slew[32] gpio_ana[39] gpio_pulldown[20]
+ gpio_oe[26] gpio_in[42] gpio_drive0[20] gpio_drive1[14] gpio_out[12] gpio[31] gpio_drive0[37]
+ gpio[34] gpio_pulldown[18] gpio_loopback_one[42] gpio[8] gpio_pullup[2] gpio_out[18]
+ gpio_schmitt[3] gpio_ie[42] gpio_out[16] gpio_pulldown[7] gpio_pullup[21] gpio_schmitt[22]
+ gpio_pulldown[40] gpio_slew[21] gpio_pulldown[17] gpio_schmitt[17] gpio_pulldown[26]
+ gpio_pulldown[35] gpio_drive1[31] gpio_slew[1] gpio_ana[17] gpio_oe[4] gpio_slew[11]
+ gpio_slew[20] gpio_slew[19] gpio_slew[40] gpio[17] gpio_oe[14] vccd gpio_drive1[40]
+ gpio_in[23] gpio_oe[23] gpio_oe[32] gpio_in[21] gpio_drive0[31] gpio[38] gpio_drive1[25]
+ gpio_pullup[43] gpio[18] gpio_loopback_one[39] gpio_pullup[23] gpio_drive0[40] gpio[5]
+ gpio_drive0[25] gpio_drive1[19] gpio_in[24] gpio_schmitt[41] gpio_schmitt[0] gpio[27]
+ gpio_pulldown[4] gpio_slew[42] gpio_schmitt[10] gpio_pulldown[14] gpio_ie[8] gpio_pulldown[23]
+ gpio[28] gpio_pulldown[32] gpio_oe[21] gpio_ie[18] gpio_ie[27] gpio_ie[36] gpio_ana[38]
+ gpio_out[38] gpio_drive0[19] gpio_drive1[4] gpio[7] gpio_oe[1] gpio[12] gpio_oe[11]
+ gpio_oe[20] gpio_oe[40] gpio_ie[22] gpio_drive1[36] gpio_pullup[16] vddio gpio_ie[39]
+ gpio[15] resetb gpio_drive0[4] gpio[37] gpio_in[41] gpio_schmitt[38] gpio_out[40]
+ vssd
Xgf180mcu_ocd_io__fill10_912 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_923 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_934 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_945 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_956 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_967 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_978 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_901 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_989 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_19 vccd gpio_loopback_one[12] gpio_loopback_zero[12] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_720 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_731 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_742 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_208 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_219 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_753 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_764 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_775 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_786 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_797 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[6] vddio gpio_drive0[6] gpio_drive1[6] gpio_pullup[6] vccd gpio_ana[6] gpio_out[6]
+ gpio_ie[6] gpio[6] gpio_slew[6] gpio_in[6] gpio_oe[6] gpio_pulldown[6] gpio_schmitt[6]
+ vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_550 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_561 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_572 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_583 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_594 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill5_2 vccd vssd vddio vssd gf180mcu_ocd_io__fill5
Xgf180mcu_ocd_io__fill10x_9 vccd gpio_loopback_one[2] gpio_loopback_zero[2] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_391 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_380 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgpio_42_pad vddio gpio_drive0[42] gpio_drive1[42] gpio_pullup[42] vccd gpio_ana[42]
+ gpio_out[42] gpio_ie[42] gpio[42] gpio_slew[42] gpio_in[42] gpio_oe[42] gpio_pulldown[42]
+ gpio_schmitt[42] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_1040 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_902 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_913 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_924 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_935 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_946 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_957 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_979 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_209 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_710 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_721 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_732 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_743 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_754 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_765 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_776 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_787 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_798 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[5] vddio gpio_drive0[5] gpio_drive1[5] gpio_pullup[5] vccd gpio_ana[5] gpio_out[5]
+ gpio_ie[5] gpio[5] gpio_slew[5] gpio_in[5] gpio_oe[5] gpio_pulldown[5] gpio_schmitt[5]
+ vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_540 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_551 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_562 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_573 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_584 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_595 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_392 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_381 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_370 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1041 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1030 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_903 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_914 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_936 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_947 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_958 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_925 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_700 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_711 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_722 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_733 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_744 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_755 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_766 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_777 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_788 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_799 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[4] vddio gpio_drive0[4] gpio_drive1[4] gpio_pullup[4] vccd gpio_ana[4] gpio_out[4]
+ gpio_ie[4] gpio[4] gpio_slew[4] gpio_in[4] gpio_oe[4] gpio_pulldown[4] gpio_schmitt[4]
+ vssd vssd gf180mcu_ocd_io__bi_a
Xuser1_vccd_pad vddio vssd vccd vssd gf180mcu_ocd_io__vdd
Xgf180mcu_ocd_io__fill10_530 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_541 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_552 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_563 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_574 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_585 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_596 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_393 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_382 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_371 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_360 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[29] vddio gpio_drive0[29] gpio_drive1[29] gpio_pullup[29] vccd gpio_ana[29]
+ gpio_out[29] gpio_ie[29] gpio[29] gpio_slew[29] gpio_in[29] gpio_oe[29] gpio_pulldown[29]
+ gpio_schmitt[29] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_190 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1042 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1031 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1020 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_904 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_926 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_937 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_948 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_959 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_701 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_712 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_723 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_734 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_745 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_756 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_767 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_778 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_789 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[3] vddio gpio_drive0[3] gpio_drive1[3] gpio_pullup[3] vccd gpio_ana[3] gpio_out[3]
+ gpio_ie[3] gpio[3] gpio_slew[3] gpio_in[3] gpio_oe[3] gpio_pulldown[3] gpio_schmitt[3]
+ vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_520 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_531 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_542 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_553 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_564 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_575 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_586 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_597 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_394 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_383 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_372 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_361 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_350 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[28] vddio gpio_drive0[28] gpio_drive1[28] gpio_pullup[28] vccd gpio_ana[28]
+ gpio_out[28] gpio_ie[28] gpio[28] gpio_slew[28] gpio_in[28] gpio_oe[28] gpio_pulldown[28]
+ gpio_schmitt[28] vssd vssd gf180mcu_ocd_io__bi_a
Xsimple_por_0 vddio porb_h por_h vssd simple_por
Xvssa_pad vddio vssd vccd vssd gf180mcu_ocd_io__dvss
Xgf180mcu_ocd_io__fill10_180 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_191 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1043 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1032 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1021 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1010 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_905 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_927 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_938 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_949 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_916 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_702 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_713 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_724 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_735 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_746 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_757 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_768 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_779 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[2] vddio gpio_drive0[2] gpio_drive1[2] gpio_pullup[2] vccd gpio_ana[2] gpio_out[2]
+ gpio_ie[2] gpio[2] gpio_slew[2] gpio_in[2] gpio_oe[2] gpio_pulldown[2] gpio_schmitt[2]
+ vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_521 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_532 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_543 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_554 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_565 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_576 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_587 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_598 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_510 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[27] vddio gpio_drive0[27] gpio_drive1[27] gpio_pullup[27] vccd gpio_ana[27]
+ gpio_out[27] gpio_ie[27] gpio[27] gpio_slew[27] gpio_in[27] gpio_oe[27] gpio_pulldown[27]
+ gpio_schmitt[27] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_395 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_384 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_373 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_362 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_351 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_340 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_181 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_192 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1044 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1033 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1022 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1011 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1000 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_906 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_917 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_928 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xvddio_pad_0 vccd vssd vddio vssd gf180mcu_ocd_io__dvdd
Xgf180mcu_ocd_io__fill10_703 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_714 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_736 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_769 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[1] vddio gpio_drive0[1] gpio_drive1[1] gpio_pullup[1] vccd gpio_ana[1] gpio_out[1]
+ gpio_ie[1] gpio[1] gpio_slew[1] gpio_in[1] gpio_oe[1] gpio_pulldown[1] gpio_schmitt[1]
+ vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_522 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_533 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_544 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_555 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_566 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_577 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_588 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_599 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_511 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_500 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[26] vddio gpio_drive0[26] gpio_drive1[26] gpio_pullup[26] vccd gpio_ana[26]
+ gpio_out[26] gpio_ie[26] gpio[26] gpio_slew[26] gpio_in[26] gpio_oe[26] gpio_pulldown[26]
+ gpio_schmitt[26] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_396 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_385 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_374 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_363 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_352 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_341 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_330 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_182 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1034 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1001 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xvddio_pad_1 vccd vssd vddio vssd gf180mcu_ocd_io__dvdd
Xgf180mcu_ocd_io__fill10_907 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_918 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_929 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xuser2_corner vccd vddio vssd gf180mcu_ocd_io__cor
Xgf180mcu_ocd_io__fill10_715 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_726 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_737 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_748 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_759 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[0] vddio gpio_drive0[0] gpio_drive1[0] gpio_pullup[0] vccd gpio_ana[0] gpio_out[0]
+ gpio_ie[0] gpio[0] gpio_slew[0] gpio_in[0] gpio_oe[0] gpio_pulldown[0] gpio_schmitt[0]
+ vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_523 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_534 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_556 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_567 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_578 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_589 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_512 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_501 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xuser2_vssa_pad vddio vssd vccd vssd gf180mcu_ocd_io__dvss
Xvssd_pad vccd vssd vddio vssd gf180mcu_ocd_io__vss
Xgf180mcu_ocd_io__fill10_397 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_386 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_375 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_364 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_353 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_342 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_320 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[25] vddio gpio_drive0[25] gpio_drive1[25] gpio_pullup[25] vccd gpio_ana[25]
+ gpio_out[25] gpio_ie[25] gpio[25] gpio_slew[25] gpio_in[25] gpio_oe[25] gpio_pulldown[25]
+ gpio_schmitt[25] vssd vssd gf180mcu_ocd_io__bi_a
Xgpio_39_pad vddio gpio_drive0[40] gpio_drive1[40] gpio_pullup[40] vccd gpio_ana[40]
+ gpio_out[40] gpio_ie[40] gpio[40] gpio_slew[40] gpio_in[40] gpio_oe[40] gpio_pulldown[40]
+ gpio_schmitt[40] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_150 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_183 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1035 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1002 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_908 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_919 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_705 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_716 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_727 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_738 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_749 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_513 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_524 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_502 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_535 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_546 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_557 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_568 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_579 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_398 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_376 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_365 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_354 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_343 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_332 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_321 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_310 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[24] vddio gpio_drive0[24] gpio_drive1[24] gpio_pullup[24] vccd gpio_ana[24]
+ gpio_out[24] gpio_ie[24] gpio[24] gpio_slew[24] gpio_in[24] gpio_oe[24] gpio_pulldown[24]
+ gpio_schmitt[24] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_140 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_151 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_184 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_195 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1036 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1025 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1014 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1003 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_909 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10y_0 vccd vssd porb_h porb_l vddio vssd gf180mcu_ocd_io__fill10y
Xgf180mcu_ocd_io__fill10_706 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_717 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_728 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_739 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_525 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_536 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_547 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_558 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_569 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_503 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_399 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_388 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_377 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_366 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_355 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_344 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_333 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_322 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_311 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_300 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[23] vddio gpio_drive0[23] gpio_drive1[23] gpio_pullup[23] vccd gpio_ana[23]
+ gpio_out[23] gpio_ie[23] gpio[23] gpio_slew[23] gpio_in[23] gpio_oe[23] gpio_pulldown[23]
+ gpio_schmitt[23] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_130 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_141 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_152 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_185 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_196 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1015 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1004 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1026 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_707 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_718 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_729 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xuser2_vssd_pad vccd vssd vddio vssd gf180mcu_ocd_io__vss
Xgf180mcu_ocd_io__fill10_526 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_515 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_537 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_548 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_559 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_504 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xvdda_pad vccd vssd vddio vssd gf180mcu_ocd_io__dvdd
Xpads[22] vddio gpio_drive0[22] gpio_drive1[22] gpio_pullup[22] vccd gpio_ana[22]
+ gpio_out[22] gpio_ie[22] gpio[22] gpio_slew[22] gpio_in[22] gpio_oe[22] gpio_pulldown[22]
+ gpio_schmitt[22] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_389 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_378 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_367 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_356 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_345 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_334 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_323 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_312 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_301 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_890 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_120 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_131 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_142 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_153 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_175 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_186 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_197 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1038 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1027 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1016 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1005 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_708 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_719 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_527 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_516 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_538 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_549 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_505 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[21] vddio gpio_drive0[21] gpio_drive1[21] gpio_pullup[21] vccd gpio_ana[21]
+ gpio_out[21] gpio_ie[21] gpio[21] gpio_slew[21] gpio_in[21] gpio_oe[21] gpio_pulldown[21]
+ gpio_schmitt[21] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_379 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_368 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_357 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_346 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_335 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_324 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_313 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_302 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_880 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_891 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_110 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_132 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_143 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_154 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_176 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_187 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_198 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1039 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1028 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1017 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1006 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_709 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_517 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_528 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_539 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_506 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_369 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_358 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_347 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_336 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_325 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_314 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[20] vddio gpio_drive0[20] gpio_drive1[20] gpio_pullup[20] vccd gpio_ana[20]
+ gpio_out[20] gpio_ie[20] gpio[20] gpio_slew[20] gpio_in[20] gpio_oe[20] gpio_pulldown[20]
+ gpio_schmitt[20] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_881 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_892 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_100 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_111 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_122 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_133 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_144 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_155 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_177 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_188 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_199 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgpio_41_pad vddio gpio_drive0[41] gpio_drive1[41] gpio_pullup[41] vccd gpio_ana[41]
+ gpio_out[41] gpio_ie[41] gpio[41] gpio_slew[41] gpio_in[41] gpio_oe[41] gpio_pulldown[41]
+ gpio_schmitt[41] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_1029 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1018 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1007 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_518 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_529 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_507 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xuser2_vdda_pad vccd vssd vddio vssd gf180mcu_ocd_io__dvdd
Xgf180mcu_ocd_io__fill10_359 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_348 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_337 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_326 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_315 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_304 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_860 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_882 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_893 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_871 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_112 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_123 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_134 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_145 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_156 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_189 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_690 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1019 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1008 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_519 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_508 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_349 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_338 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_327 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_316 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_305 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_850 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_861 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_872 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_883 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_894 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_102 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_113 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_124 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_135 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_146 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_157 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_179 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_680 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_691 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1009 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_509 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_306 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_840 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_851 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_862 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_339 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_328 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_873 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_884 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_895 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_103 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_114 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_125 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_136 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_147 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_670 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_681 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_692 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_90 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_329 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_318 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_307 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10z_10 vddio vssd vccd vssd mask_rev[20] mask_rev[21] gf180mcu_ocd_io__fill10z
Xgf180mcu_ocd_io__fill10_830 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_852 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_863 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_874 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_896 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_104 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_115 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_126 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_137 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_148 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_660 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_671 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_682 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_693 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xuser_id_programming_0 mask_rev[0] mask_rev[10] mask_rev[11] mask_rev[12] mask_rev[13]
+ mask_rev[14] mask_rev[15] mask_rev[16] mask_rev[17] mask_rev[18] mask_rev[19] mask_rev[1]
+ mask_rev[20] mask_rev[21] mask_rev[22] mask_rev[23] mask_rev[24] mask_rev[25] mask_rev[26]
+ mask_rev[27] mask_rev[28] mask_rev[29] mask_rev[2] mask_rev[30] mask_rev[31] mask_rev[3]
+ mask_rev[4] mask_rev[5] mask_rev[6] mask_rev[7] mask_rev[8] mask_rev[9] vccd vssd
+ user_id_programming
Xgf180mcu_ocd_io__fill10_490 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_80 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_91 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_319 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_308 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_820 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_831 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_842 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_853 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_864 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_875 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_897 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10z_11 vddio vssd vccd vssd mask_rev[22] mask_rev[23] gf180mcu_ocd_io__fill10z
Xgf180mcu_ocd_io__fill10_886 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_105 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_116 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_127 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_149 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_650 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_661 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_672 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_683 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_694 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_491 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_480 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_81 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_70 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_92 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_309 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_810 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_821 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_832 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_843 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_854 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_865 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_876 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_887 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_898 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10z_12 vddio vssd vccd vssd mask_rev[24] mask_rev[25] gf180mcu_ocd_io__fill10z
Xgpio_38_pad vddio gpio_drive0[39] gpio_drive1[39] gpio_pullup[39] vccd gpio_ana[39]
+ gpio_out[39] gpio_ie[39] gpio[39] gpio_slew[39] gpio_in[39] gpio_oe[39] gpio_pulldown[39]
+ gpio_schmitt[39] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_106 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_117 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_128 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_139 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_640 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_651 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_662 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_673 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_684 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_695 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_492 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_481 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_470 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xresetb_pad vddio resetb_pulldown resetb_pullup vccd resetb resetb_core vssd vssd
+ gf180mcu_ocd_io__in_s
Xgf180mcu_ocd_io__fill10_82 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_71 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_60 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_93 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_0 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_811 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_822 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_833 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_844 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_866 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_877 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_888 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_899 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10z_13 vddio vssd vccd vssd mask_rev[26] mask_rev[27] gf180mcu_ocd_io__fill10z
Xgf180mcu_ocd_io__fill10_800 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_107 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_118 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_129 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_630 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_641 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_652 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_663 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_674 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_685 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_696 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_493 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_482 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_471 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_460 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_290 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_83 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_72 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_61 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_50 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_94 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_1 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_801 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_812 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_823 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_834 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_845 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_867 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10z_14 vddio vssd vccd vssd mask_rev[28] mask_rev[29] gf180mcu_ocd_io__fill10z
Xgf180mcu_ocd_io__fill10_856 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_878 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_889 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_108 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_119 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_620 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_631 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_642 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_653 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_664 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_675 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_686 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_697 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_494 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_483 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_472 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_461 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_450 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xuser1_vssd_pad vccd vssd vddio vssd gf180mcu_ocd_io__vss
Xgf180mcu_ocd_io__fill10_291 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_95 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_84 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_73 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_62 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_51 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_40 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_280 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_2 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10z_15 vddio vssd vccd vssd mask_rev[30] mask_rev[31] gf180mcu_ocd_io__fill10z
Xgf180mcu_ocd_io__fill10_802 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_813 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_824 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_835 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_846 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_857 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_868 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_879 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_109 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_610 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_621 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_632 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_643 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_654 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_665 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_676 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_687 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_698 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_495 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_484 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_473 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_462 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_451 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_440 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[37] vddio gpio_drive0[37] gpio_drive1[37] gpio_pullup[37] vccd gpio_ana[37]
+ gpio_out[37] gpio_ie[37] gpio[37] gpio_slew[37] gpio_in[37] gpio_oe[37] gpio_pulldown[37]
+ gpio_schmitt[37] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_292 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_96 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_85 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_74 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_63 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_52 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_41 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_30 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_270 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_281 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_3 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_803 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_814 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_825 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_836 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_858 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_869 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10z_16 vddio vssd vccd vssd por_h porb_h gf180mcu_ocd_io__fill10z
Xgf180mcu_ocd_io__fill10_847 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_600 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_611 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_622 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_633 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_644 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_655 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_677 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_688 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_699 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_496 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_474 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_463 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_452 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_441 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_430 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[36] vddio gpio_drive0[36] gpio_drive1[36] gpio_pullup[36] vccd gpio_ana[36]
+ gpio_out[36] gpio_ie[36] gpio[36] gpio_slew[36] gpio_in[36] gpio_oe[36] gpio_pulldown[36]
+ gpio_schmitt[36] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_293 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_86 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_97 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_75 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_64 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_53 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_42 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_31 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_20 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_271 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_282 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[19] vddio gpio_drive0[19] gpio_drive1[19] gpio_pullup[19] vccd gpio_ana[19]
+ gpio_out[19] gpio_ie[19] gpio[19] gpio_slew[19] gpio_in[19] gpio_oe[19] gpio_pulldown[19]
+ gpio_schmitt[19] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_4 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_804 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_815 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_826 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_837 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_848 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_859 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_601 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_612 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_623 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_634 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_645 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_656 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_667 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_678 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_497 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_486 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_475 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_464 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_453 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_442 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_431 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_420 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[35] vddio gpio_drive0[35] gpio_drive1[35] gpio_pullup[35] vccd gpio_ana[35]
+ gpio_out[35] gpio_ie[35] gpio[35] gpio_slew[35] gpio_in[35] gpio_oe[35] gpio_pulldown[35]
+ gpio_schmitt[35] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_294 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_87 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_65 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_76 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_54 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_43 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_32 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_21 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_10 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_98 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_250 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_272 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_283 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[18] vddio gpio_drive0[18] gpio_drive1[18] gpio_pullup[18] vccd gpio_ana[18]
+ gpio_out[18] gpio_ie[18] gpio[18] gpio_slew[18] gpio_in[18] gpio_oe[18] gpio_pulldown[18]
+ gpio_schmitt[18] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_5 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_805 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_816 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_838 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_849 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_827 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_602 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_613 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_624 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_635 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_646 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_657 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_668 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_679 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_498 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_487 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_476 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_465 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_454 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_432 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_421 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_410 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[34] vddio gpio_drive0[34] gpio_drive1[34] gpio_pullup[34] vccd gpio_ana[34]
+ gpio_out[34] gpio_ie[34] gpio[34] gpio_slew[34] gpio_in[34] gpio_oe[34] gpio_pulldown[34]
+ gpio_schmitt[34] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10x_40 vccd gpio_loopback_one[33] gpio_loopback_zero[33] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_295 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_240 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_251 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_262 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_273 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_284 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[17] vddio gpio_drive0[17] gpio_drive1[17] gpio_pullup[17] vccd gpio_ana[17]
+ gpio_out[17] gpio_ie[17] gpio[17] gpio_slew[17] gpio_in[17] gpio_oe[17] gpio_pulldown[17]
+ gpio_schmitt[17] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_66 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_77 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_44 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_55 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_33 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_22 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_11 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_88 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_99 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10z_0 vddio vssd vccd vssd mask_rev[0] mask_rev[1] gf180mcu_ocd_io__fill10z
Xgf180mcu_ocd_io__fill10_6 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_806 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_817 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_839 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_603 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_614 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_625 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_636 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_647 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_658 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_669 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xvccd_pad vddio vssd vccd vssd gf180mcu_ocd_io__vdd
Xgf180mcu_ocd_io__fill10_499 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_488 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_477 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_466 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_455 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_444 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_433 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_422 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_411 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_400 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[33] vddio gpio_drive0[33] gpio_drive1[33] gpio_pullup[33] vccd gpio_ana[33]
+ gpio_out[33] gpio_ie[33] gpio[33] gpio_slew[33] gpio_in[33] gpio_oe[33] gpio_pulldown[33]
+ gpio_schmitt[33] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10x_30 vccd gpio_loopback_one[23] gpio_loopback_zero[23] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_41 vccd gpio_loopback_one[34] gpio_loopback_zero[34] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_230 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_241 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_252 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_263 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_274 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[16] vddio gpio_drive0[16] gpio_drive1[16] gpio_pullup[16] vccd gpio_ana[16]
+ gpio_out[16] gpio_ie[16] gpio[16] gpio_slew[16] gpio_in[16] gpio_oe[16] gpio_pulldown[16]
+ gpio_schmitt[16] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_296 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_285 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_67 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_45 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_56 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_34 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_23 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_12 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_78 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_89 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10z_1 vddio vssd vccd vssd mask_rev[2] mask_rev[3] gf180mcu_ocd_io__fill10z
Xgf180mcu_ocd_io__fill10_7 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_807 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_829 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__bi_a_0 vddio gpio_drive0[38] gpio_drive2[38] gpio_pullup[38] vccd
+ gpio_ana[38] gpio_out[38] gpio_ie[38] gpio[38] gpio_slew[38] gpio_in[38] gpio_oe[38]
+ gpio_pulldown[38] gpio_schmitt[38] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_818 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_604 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_615 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_626 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_637 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_648 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_659 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgpio_43_pad vddio gpio_drive0[43] gpio_drive1[43] gpio_pullup[43] vccd gpio_ana[43]
+ gpio_out[43] gpio_ie[43] gpio[43] gpio_slew[43] gpio_in[43] gpio_oe[43] gpio_pulldown[43]
+ gpio_schmitt[43] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_489 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_478 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_467 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_456 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_445 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_434 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_423 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_412 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[32] vddio gpio_drive0[32] gpio_drive1[32] gpio_pullup[32] vccd gpio_ana[32]
+ gpio_out[32] gpio_ie[32] gpio[32] gpio_slew[32] gpio_in[32] gpio_oe[32] gpio_pulldown[32]
+ gpio_schmitt[32] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_990 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_31 vccd gpio_loopback_one[24] gpio_loopback_zero[24] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_20 vccd gpio_loopback_one[13] gpio_loopback_zero[13] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xpads[15] vddio gpio_drive0[15] gpio_drive1[15] gpio_pullup[15] vccd gpio_ana[15]
+ gpio_out[15] gpio_ie[15] gpio[15] gpio_slew[15] gpio_in[15] gpio_oe[15] gpio_pulldown[15]
+ gpio_schmitt[15] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_297 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_79 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_68 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_46 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_57 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_35 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_24 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_13 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_220 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_231 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_242 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_253 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_264 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_286 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_42 vccd gpio_loopback_one[35] gpio_loopback_zero[35] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10z_2 vddio vssd vccd vssd mask_rev[4] mask_rev[5] gf180mcu_ocd_io__fill10z
Xgf180mcu_ocd_io__fill10_8 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_808 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_819 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_605 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_616 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_627 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_638 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_649 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_479 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_468 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_446 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_435 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_424 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_413 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_402 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[31] vddio gpio_drive0[31] gpio_drive1[31] gpio_pullup[31] vccd gpio_ana[31]
+ gpio_out[31] gpio_ie[31] gpio[31] gpio_slew[31] gpio_in[31] gpio_oe[31] gpio_pulldown[31]
+ gpio_schmitt[31] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_980 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_991 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_21 vccd gpio_loopback_one[14] gpio_loopback_zero[14] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xpads[14] vddio gpio_drive0[14] gpio_drive1[14] gpio_pullup[14] vccd gpio_ana[14]
+ gpio_out[14] gpio_ie[14] gpio[14] gpio_slew[14] gpio_in[14] gpio_oe[14] gpio_pulldown[14]
+ gpio_schmitt[14] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10x_32 vccd gpio_loopback_one[25] gpio_loopback_zero[25] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_298 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_10 vccd gpio_loopback_one[3] gpio_loopback_zero[3] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_287 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_69 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_58 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_47 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_36 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_25 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_14 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_210 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_221 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_232 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_243 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_254 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_43 vccd gpio_loopback_one[36] gpio_loopback_zero[36] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_265 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_276 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10z_3 vddio vssd vccd vssd mask_rev[6] mask_rev[7] gf180mcu_ocd_io__fill10z
Xgf180mcu_ocd_io__fill10_9 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xuser2_vccd_pad vddio vssd vccd vssd gf180mcu_ocd_io__vdd
Xgf180mcu_ocd_io__fill10x_0 vccd resetb_loopback_one resetb_loopback_zero vddio vssd
+ vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_809 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_617 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_639 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_469 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_458 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_447 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_436 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_425 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_414 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_403 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xuser1_vssa_pad_0 vddio vssd vccd vssd gf180mcu_ocd_io__dvss
Xpads[30] vddio gpio_drive0[30] gpio_drive1[30] gpio_pullup[30] vccd gpio_ana[30]
+ gpio_out[30] gpio_ie[30] gpio[30] gpio_slew[30] gpio_in[30] gpio_oe[30] gpio_pulldown[30]
+ gpio_schmitt[30] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_970 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_981 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_992 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_22 vccd gpio_loopback_one[15] gpio_loopback_zero[15] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_33 vccd gpio_loopback_one[26] gpio_loopback_zero[26] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_11 vccd gpio_loopback_one[4] gpio_loopback_zero[4] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_299 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_288 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_48 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_26 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_15 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_200 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_211 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_222 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_233 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_244 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_255 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_44 vccd gpio_loopback_one[37] gpio_loopback_zero[37] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_266 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_277 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[13] vddio gpio_drive0[13] gpio_drive1[13] gpio_pullup[13] vccd gpio_ana[13]
+ gpio_out[13] gpio_ie[13] gpio[13] gpio_slew[13] gpio_in[13] gpio_oe[13] gpio_pulldown[13]
+ gpio_schmitt[13] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10z_4 vddio vssd vccd vssd mask_rev[8] mask_rev[9] gf180mcu_ocd_io__fill10z
Xgf180mcu_ocd_io__fill10x_1 vccd gpio_loopback_one[38] gpio_loopback_zero[38] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_607 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_618 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_629 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_404 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_459 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_448 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_437 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_426 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_960 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_971 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xuser1_vssa_pad_1 vddio vssd vccd vssd gf180mcu_ocd_io__dvss
Xgf180mcu_ocd_io__fill10_982 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_993 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_23 vccd gpio_loopback_one[16] gpio_loopback_zero[16] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_34 vccd gpio_loopback_one[27] gpio_loopback_zero[27] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_12 vccd gpio_loopback_one[5] gpio_loopback_zero[5] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_201 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_212 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_223 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_234 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_245 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_256 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_267 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_278 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_790 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[12] vddio gpio_drive0[12] gpio_drive1[12] gpio_pullup[12] vccd gpio_ana[12]
+ gpio_out[12] gpio_ie[12] gpio[12] gpio_slew[12] gpio_in[12] gpio_oe[12] gpio_pulldown[12]
+ gpio_schmitt[12] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_49 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_27 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_16 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xvssio_pad_0 vddio vssd vccd vssd gf180mcu_ocd_io__dvss
Xgf180mcu_ocd_io__fill10z_5 vddio vssd vccd vssd mask_rev[10] mask_rev[11] gf180mcu_ocd_io__fill10z
Xgf180mcu_ocd_io__fill10x_2 vccd gpio_loopback_one[39] gpio_loopback_zero[39] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_608 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_619 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_449 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_438 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_427 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_416 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_405 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_950 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_961 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_972 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_994 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_24 vccd gpio_loopback_one[17] gpio_loopback_zero[17] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_35 vccd gpio_loopback_one[28] gpio_loopback_zero[28] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_13 vccd gpio_loopback_one[6] gpio_loopback_zero[6] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_202 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_213 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_224 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_246 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_257 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_268 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_279 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_780 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_791 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[11] vddio gpio_drive0[11] gpio_drive1[11] gpio_pullup[11] vccd gpio_ana[11]
+ gpio_out[11] gpio_ie[11] gpio[11] gpio_slew[11] gpio_in[11] gpio_oe[11] gpio_pulldown[11]
+ gpio_schmitt[11] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_39 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_28 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_17 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xvssio_pad_1 vddio vssd vccd vssd gf180mcu_ocd_io__dvss
Xgf180mcu_ocd_io__fill10z_6 vddio vssd vccd vssd mask_rev[12] mask_rev[13] gf180mcu_ocd_io__fill10z
Xgf180mcu_ocd_io__fill10x_3 vccd gpio_loopback_one[40] gpio_loopback_zero[40] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_609 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_439 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_428 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_417 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_406 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_940 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_951 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_962 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_973 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_995 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_25 vccd gpio_loopback_one[18] gpio_loopback_zero[18] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_36 vccd gpio_loopback_one[29] gpio_loopback_zero[29] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_14 vccd gpio_loopback_one[7] gpio_loopback_zero[7] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xpads[10] vddio gpio_drive0[10] gpio_drive1[10] gpio_pullup[10] vccd gpio_ana[10]
+ gpio_out[10] gpio_ie[10] gpio[10] gpio_slew[10] gpio_in[10] gpio_oe[10] gpio_pulldown[10]
+ gpio_schmitt[10] vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10_29 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_18 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_203 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_214 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_225 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_247 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_258 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_269 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_770 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_781 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_792 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10z_7 vddio vssd vccd vssd mask_rev[14] mask_rev[15] gf180mcu_ocd_io__fill10z
Xgf180mcu_ocd_io__fill10x_4 vccd gpio_loopback_one[41] gpio_loopback_zero[41] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_418 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_407 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_930 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_941 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_952 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_963 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_974 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_985 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xcorner[1] vccd vddio vssd gf180mcu_ocd_io__cor
Xgf180mcu_ocd_io__fill10_996 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_26 vccd gpio_loopback_one[19] gpio_loopback_zero[19] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_15 vccd gpio_loopback_one[8] gpio_loopback_zero[8] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_37 vccd gpio_loopback_one[30] gpio_loopback_zero[30] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_19 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_204 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_215 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_226 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_259 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_248 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_760 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_771 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_782 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_793 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_590 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10z_8 vddio vssd vccd vssd mask_rev[16] mask_rev[17] gf180mcu_ocd_io__fill10z
Xgf180mcu_ocd_io__fill10x_5 vccd gpio_loopback_one[42] gpio_loopback_zero[42] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_419 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_408 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_920 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_931 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_942 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_964 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_975 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xcorner[0] vccd vddio vssd gf180mcu_ocd_io__cor
Xgf180mcu_ocd_io__fill10_986 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_27 vccd gpio_loopback_one[20] gpio_loopback_zero[20] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_16 vccd gpio_loopback_one[9] gpio_loopback_zero[9] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_38 vccd gpio_loopback_one[31] gpio_loopback_zero[31] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_205 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_216 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_227 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_238 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_249 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_750 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_783 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_794 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_761 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[9] vddio gpio_drive0[9] gpio_drive1[9] gpio_pullup[9] vccd gpio_ana[9] gpio_out[9]
+ gpio_ie[9] gpio[9] gpio_slew[9] gpio_in[9] gpio_oe[9] gpio_pulldown[9] gpio_schmitt[9]
+ vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill10z_9 vddio vssd vccd vssd mask_rev[18] mask_rev[19] gf180mcu_ocd_io__fill10z
Xgf180mcu_ocd_io__fill10_580 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_591 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_6 vccd gpio_loopback_one[43] gpio_loopback_zero[43] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xuser1_vdda_pad_0 vccd vssd vddio vssd gf180mcu_ocd_io__dvdd
Xgf180mcu_ocd_io__fill10_409 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_910 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_921 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_932 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_943 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_965 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_976 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_987 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_28 vccd gpio_loopback_one[21] gpio_loopback_zero[21] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_17 vccd gpio_loopback_one[10] gpio_loopback_zero[10] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_39 vccd gpio_loopback_one[32] gpio_loopback_zero[32] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_206 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_217 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_228 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_239 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_740 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_751 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_762 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_784 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_795 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_773 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[8] vddio gpio_drive0[8] gpio_drive1[8] gpio_pullup[8] vccd gpio_ana[8] gpio_out[8]
+ gpio_ie[8] gpio[8] gpio_slew[8] gpio_in[8] gpio_oe[8] gpio_pulldown[8] gpio_schmitt[8]
+ vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill5_0 vccd vssd vddio vssd gf180mcu_ocd_io__fill5
Xgf180mcu_ocd_io__fill10_570 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_581 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_592 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_7 vccd gpio_loopback_one[0] gpio_loopback_zero[0] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xuser1_vdda_pad_1 vccd vssd vddio vssd gf180mcu_ocd_io__dvdd
Xgf180mcu_ocd_io__fill10_911 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_922 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_933 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_944 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_955 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_966 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_977 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_988 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_999 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_29 vccd gpio_loopback_one[22] gpio_loopback_zero[22] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10x_18 vccd gpio_loopback_one[11] gpio_loopback_zero[11] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xgf180mcu_ocd_io__fill10_207 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_218 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_229 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_730 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_741 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_752 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_763 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_774 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_796 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_785 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xpads[7] vddio gpio_drive0[7] gpio_drive1[7] gpio_pullup[7] vccd gpio_ana[7] gpio_out[7]
+ gpio_ie[7] gpio[7] gpio_slew[7] gpio_in[7] gpio_oe[7] gpio_pulldown[7] gpio_schmitt[7]
+ vssd vssd gf180mcu_ocd_io__bi_a
Xgf180mcu_ocd_io__fill5_1 vccd vssd vddio vssd gf180mcu_ocd_io__fill5
Xgf180mcu_ocd_io__fill10_560 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_571 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10_593 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
Xgf180mcu_ocd_io__fill10x_8 vccd gpio_loopback_one[1] gpio_loopback_zero[1] vddio
+ vssd vssd gf180mcu_ocd_io__fill10x
Xuser1_corner vccd vddio vssd gf180mcu_ocd_io__cor
Xgf180mcu_ocd_io__fill10_390 vccd vssd vddio vssd gf180mcu_ocd_io__fill10
.ends

.subckt horz_connects_gpio_disabled m1_0_133# m1_1576_37# m2_15068_0# m1_932_37# m1_1074_37#
+ m1_13244_37# m1_182_37# m1_703_37# m1_13390_36# m1_1787_37# m1_13536_37#
X0 m1_0_133# m1_932_37# rm1 r_width=0.38u r_length=85n
X1 m1_0_133# m1_1074_37# rm1 r_width=0.38u r_length=85n
X2 m1_0_133# m1_703_37# rm1 r_width=0.38u r_length=85n
X3 m1_0_133# m1_13244_37# rm1 r_width=0.38u r_length=85n
X4 m1_0_133# m1_13536_37# rm1 r_width=0.38u r_length=85n
X5 m1_0_133# m1_1787_37# rm1 r_width=0.38u r_length=85n
X6 m1_0_133# m1_1576_37# rm1 r_width=0.38u r_length=85n
X7 m1_0_133# m1_182_37# rm1 r_width=0.38u r_length=85n
X8 m1_0_133# m1_13390_36# rm1 r_width=0.38u r_length=85n
.ends

.subckt vert_connects_gpio_disabled m3_0_120# m3_0_14444# m3_0_13800# m3_0_15194#
+ m2_32_14673# m3_0_14302# m2_32_14444# m2_32_13800# m2_32_15194# m2_32_14302# m3_0_1840#
+ m3_0_1986# m2_32_1840# m2_32_1986# m3_0_308# m3_0_2132# m2_32_2132# m3_0_13589#
+ m2_32_13589# m3_0_14673#
X0 m3_0_15194# m3_0_120# rm4 r_width=0.38u r_length=80n
X1 m3_0_14302# m3_0_120# rm4 r_width=0.38u r_length=80n
X2 m3_0_14444# m3_0_120# rm4 r_width=0.38u r_length=80n
X3 m3_0_13589# m3_0_120# rm4 r_width=0.38u r_length=80n
X4 m3_0_13800# m3_0_120# rm4 r_width=0.38u r_length=80n
X5 m3_0_14673# m3_0_120# rm4 r_width=0.38u r_length=80n
X6 m3_0_1986# m3_0_120# rm4 r_width=0.38u r_length=80n
X7 m3_0_1840# m3_0_120# rm4 r_width=0.38u r_length=80n
X8 m3_0_2132# m3_0_120# rm4 r_width=0.38u r_length=80n
.ends

.subckt openframe_user_project gpio_in[38] gpio_in[40] gpio_oe[40] gpio_in[39] gpio_oe[39]
+ gpio_in[41] gpio_out[41] gpio_ie[41] gpio_oe[41] gpio_in[42] gpio_out[42] gpio_ie[42]
+ gpio_oe[42] gpio_drive0[38] gpio_drive1[38] gpio_in[43] gpio_ie[38] gpio_out[38]
+ gpio_oe[38] gpio_pulldown[38] gpio_pullup[38] gpio_schmitt[38] gpio_slew[38] gpio_schmitt[42]
+ gpio_pullup[42] gpio_drive0[42] gpio_drive1[42] gpio_pulldown[42] gpio_slew[42]
+ gpio_schmitt[41] gpio_pullup[41] gpio_drive0[41] gpio_drive1[41] gpio_pulldown[41]
+ gpio_slew[41] gpio_schmitt[40] gpio_pullup[40] gpio_drive0[40] gpio_drive1[40] gpio_pulldown[40]
+ gpio_ie[40] gpio_slew[40] gpio_out[40] gpio_schmitt[39] gpio_pullup[39] gpio_drive0[39]
+ gpio_drive1[39] gpio_pulldown[39] gpio_ie[39] gpio_slew[39] gpio_out[39] gpio_out[43]
+ gpio_slew[43] gpio_ie[43] gpio_pulldown[43] gpio_drive1[43] gpio_drive0[43] gpio_pullup[43]
+ gpio_schmitt[43] gpio_oe[43] gpio_drive0[30] gpio_drive0[0] gpio_drive0[5] gpio_drive1[5]
+ gpio_drive0[6] gpio_drive1[6] gpio_drive0[7] gpio_drive1[7] gpio_drive0[8] gpio_drive1[8]
+ gpio_drive0[9] gpio_drive1[9] gpio_drive1[0] gpio_drive0[10] gpio_drive1[10] gpio_drive0[11]
+ gpio_drive1[11] gpio_drive0[12] gpio_drive1[12] gpio_drive0[13] gpio_drive1[13]
+ gpio_drive0[14] gpio_drive1[14] gpio_drive0[1] gpio_drive0[15] gpio_drive0[16] gpio_drive1[16]
+ gpio_drive0[17] gpio_drive1[17] gpio_drive0[18] gpio_drive1[18] gpio_drive0[19]
+ gpio_drive1[19] gpio_drive1[1] gpio_drive0[20] gpio_drive1[20] gpio_drive0[21] gpio_drive1[21]
+ gpio_drive0[22] gpio_drive1[22] gpio_drive0[23] gpio_drive1[23] gpio_drive0[24]
+ gpio_drive1[24] gpio_drive0[2] gpio_drive1[25] gpio_drive0[25] gpio_drive0[26] gpio_drive1[26]
+ gpio_drive0[27] gpio_drive1[27] gpio_drive0[28] gpio_drive1[28] gpio_drive0[29]
+ gpio_drive1[29] gpio_drive1[2] gpio_drive1[30] gpio_drive0[31] gpio_drive1[31] gpio_drive0[32]
+ gpio_drive1[32] gpio_drive0[33] gpio_drive1[33] gpio_drive0[34] gpio_drive1[34]
+ gpio_drive0[3] gpio_drive0[35] gpio_drive1[35] gpio_drive0[36] gpio_drive1[36] gpio_drive0[37]
+ gpio_drive1[37] gpio_drive1[3] gpio_drive0[4] gpio_drive1[4] gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[34] gpio_in[35] gpio_in[36]
+ gpio_in[37] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_ie[0] gpio_ie[10] gpio_ie[11] gpio_ie[12] gpio_ie[13] gpio_ie[14] gpio_ie[15]
+ gpio_ie[16] gpio_ie[17] gpio_ie[18] gpio_ie[19] gpio_ie[1] gpio_ie[20] gpio_ie[21]
+ gpio_ie[22] gpio_ie[23] gpio_ie[24] gpio_ie[25] gpio_ie[26] gpio_ie[27] gpio_ie[28]
+ gpio_ie[29] gpio_ie[2] gpio_ie[30] gpio_ie[31] gpio_ie[32] gpio_ie[33] gpio_ie[34]
+ gpio_ie[35] gpio_ie[36] gpio_ie[37] gpio_ie[3] gpio_ie[4] gpio_ie[5] gpio_ie[6]
+ gpio_ie[7] gpio_ie[8] gpio_ie[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[34] gpio_out[35] gpio_out[36] gpio_out[37] gpio_out[3]
+ gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] gpio_oe[0]
+ gpio_oe[10] gpio_oe[11] gpio_oe[12] gpio_oe[13] gpio_oe[14] gpio_oe[15] gpio_oe[16]
+ gpio_oe[17] gpio_oe[18] gpio_oe[19] gpio_oe[1] gpio_oe[20] gpio_oe[21] gpio_oe[22]
+ gpio_oe[23] gpio_oe[24] gpio_oe[25] gpio_oe[26] gpio_oe[27] gpio_oe[28] gpio_oe[29]
+ gpio_oe[2] gpio_oe[30] gpio_oe[31] gpio_oe[32] gpio_oe[33] gpio_oe[34] gpio_oe[35]
+ gpio_oe[36] gpio_oe[37] gpio_oe[3] gpio_oe[4] gpio_oe[5] gpio_oe[6] gpio_oe[7] gpio_oe[8]
+ gpio_oe[9] gpio_pulldown[0] gpio_pulldown[10] gpio_pulldown[11] gpio_pulldown[12]
+ gpio_pulldown[13] gpio_pulldown[14] gpio_pulldown[15] gpio_pulldown[16] gpio_pulldown[17]
+ gpio_pulldown[18] gpio_pulldown[19] gpio_pulldown[1] gpio_pulldown[20] gpio_pulldown[21]
+ gpio_pulldown[22] gpio_pulldown[23] gpio_pulldown[24] gpio_pulldown[25] gpio_pulldown[26]
+ gpio_pulldown[27] gpio_pulldown[28] gpio_pulldown[29] gpio_pulldown[2] gpio_pulldown[30]
+ gpio_pulldown[31] gpio_pulldown[32] gpio_pulldown[33] gpio_pulldown[34] gpio_pulldown[35]
+ gpio_pulldown[36] gpio_pulldown[37] gpio_pulldown[3] gpio_pulldown[4] gpio_pulldown[5]
+ gpio_pulldown[6] gpio_pulldown[7] gpio_pulldown[8] gpio_pulldown[9] gpio_pullup[0]
+ gpio_pullup[10] gpio_pullup[11] gpio_pullup[12] gpio_pullup[13] gpio_pullup[14]
+ gpio_pullup[15] gpio_pullup[16] gpio_pullup[17] gpio_pullup[18] gpio_pullup[19]
+ gpio_pullup[1] gpio_pullup[20] gpio_pullup[21] gpio_pullup[22] gpio_pullup[23] gpio_pullup[24]
+ gpio_pullup[25] gpio_pullup[26] gpio_pullup[27] gpio_pullup[28] gpio_pullup[29]
+ gpio_pullup[2] gpio_pullup[30] gpio_pullup[31] gpio_pullup[32] gpio_pullup[33] gpio_pullup[34]
+ gpio_pullup[35] gpio_pullup[36] gpio_pullup[37] gpio_pullup[3] gpio_pullup[4] gpio_pullup[5]
+ gpio_pullup[6] gpio_pullup[7] gpio_pullup[8] gpio_pullup[9] gpio_schmitt[0] gpio_schmitt[10]
+ gpio_schmitt[11] gpio_schmitt[12] gpio_schmitt[13] gpio_schmitt[14] gpio_schmitt[15]
+ gpio_schmitt[16] gpio_schmitt[17] gpio_schmitt[18] gpio_schmitt[19] gpio_schmitt[1]
+ gpio_schmitt[20] gpio_schmitt[21] gpio_schmitt[22] gpio_schmitt[23] gpio_schmitt[24]
+ gpio_schmitt[25] gpio_schmitt[26] gpio_schmitt[27] gpio_schmitt[28] gpio_schmitt[29]
+ gpio_schmitt[2] gpio_schmitt[30] gpio_schmitt[31] gpio_schmitt[32] gpio_schmitt[33]
+ gpio_schmitt[34] gpio_schmitt[35] gpio_schmitt[36] gpio_schmitt[37] gpio_schmitt[3]
+ gpio_schmitt[4] gpio_schmitt[5] gpio_schmitt[6] gpio_schmitt[7] gpio_schmitt[8]
+ gpio_schmitt[9] gpio_slew[0] gpio_slew[10] gpio_slew[11] gpio_slew[12] gpio_slew[13]
+ gpio_slew[14] gpio_slew[15] gpio_slew[16] gpio_slew[17] gpio_slew[18] gpio_slew[19]
+ gpio_slew[1] gpio_slew[20] gpio_slew[21] gpio_slew[22] gpio_slew[23] gpio_slew[24]
+ gpio_slew[25] gpio_slew[26] gpio_slew[27] gpio_slew[28] gpio_slew[29] gpio_slew[2]
+ gpio_slew[30] gpio_slew[31] gpio_slew[32] gpio_slew[33] gpio_slew[34] gpio_slew[35]
+ gpio_slew[36] gpio_slew[37] gpio_slew[3] gpio_slew[4] gpio_slew[5] gpio_slew[6]
+ gpio_slew[7] gpio_slew[8] gpio_slew[9] resetb_core gpio_ana[0] gpio_ana[1] gpio_ana[2]
+ gpio_ana[3] gpio_ana[4] gpio_ana[5] gpio_ana[6] gpio_ana[7] gpio_ana[8] gpio_ana[9]
+ gpio_ana[10] gpio_ana[11] gpio_ana[12] gpio_ana[13] gpio_ana[14] gpio_ana[15] gpio_ana[16]
+ gpio_ana[17] gpio_ana[18] gpio_ana[19] gpio_ana[20] gpio_ana[21] gpio_ana[22] gpio_ana[23]
+ gpio_ana[24] gpio_ana[25] gpio_ana[26] gpio_ana[27] gpio_ana[28] gpio_ana[29] gpio_ana[30]
+ gpio_ana[31] gpio_ana[32] gpio_ana[33] gpio_ana[34] gpio_ana[35] gpio_ana[36] gpio_ana[37]
+ gpio_ana[38] gpio_ana[39] gpio_ana[40] gpio_ana[41] gpio_ana[42] gpio_ana[43] gpio_loopback_zero[0]
+ gpio_loopback_one[0] gpio_loopback_zero[1] gpio_loopback_one[1] gpio_loopback_zero[2]
+ gpio_loopback_one[2] gpio_loopback_one[3] gpio_loopback_zero[3] gpio_loopback_zero[4]
+ gpio_loopback_one[4] gpio_loopback_one[5] gpio_loopback_zero[5] gpio_loopback_zero[6]
+ gpio_loopback_one[6] gpio_loopback_one[7] gpio_loopback_zero[7] gpio_loopback_zero[8]
+ gpio_loopback_one[8] gpio_loopback_one[9] gpio_loopback_zero[9] gpio_loopback_zero[10]
+ gpio_loopback_one[10] gpio_loopback_one[11] gpio_loopback_zero[11] gpio_loopback_zero[12]
+ gpio_loopback_one[12] gpio_loopback_one[13] gpio_loopback_zero[13] gpio_loopback_zero[14]
+ gpio_loopback_one[14] gpio_loopback_one[15] gpio_loopback_zero[15] gpio_loopback_zero[16]
+ gpio_loopback_one[16] gpio_loopback_one[17] gpio_loopback_zero[17] gpio_loopback_zero[18]
+ gpio_loopback_one[18] gpio_loopback_one[19] gpio_loopback_zero[19] gpio_loopback_zero[20]
+ gpio_loopback_one[20] gpio_loopback_one[21] gpio_loopback_zero[21] gpio_loopback_zero[22]
+ gpio_loopback_one[22] gpio_loopback_one[23] gpio_loopback_zero[23] gpio_loopback_zero[24]
+ gpio_loopback_one[24] gpio_loopback_one[25] gpio_loopback_zero[25] gpio_loopback_zero[26]
+ gpio_loopback_one[26] gpio_loopback_one[27] gpio_loopback_zero[27] gpio_loopback_zero[28]
+ gpio_loopback_one[28] gpio_loopback_one[29] gpio_loopback_zero[29] gpio_loopback_zero[30]
+ gpio_loopback_one[30] gpio_loopback_one[31] gpio_loopback_zero[31] gpio_loopback_zero[32]
+ gpio_loopback_one[32] gpio_loopback_one[33] gpio_loopback_zero[33] gpio_loopback_zero[34]
+ gpio_loopback_one[34] gpio_loopback_one[35] gpio_loopback_zero[35] gpio_loopback_zero[36]
+ gpio_loopback_one[36] gpio_loopback_one[37] gpio_loopback_zero[37] gpio_loopback_zero[38]
+ gpio_loopback_one[38] gpio_loopback_one[39] gpio_loopback_zero[39] gpio_loopback_zero[40]
+ gpio_loopback_one[40] gpio_loopback_one[41] gpio_loopback_zero[41] gpio_loopback_zero[42]
+ gpio_loopback_one[42] gpio_loopback_one[43] gpio_loopback_zero[43] resetb_pullup
+ resetb_pulldown resetb_loopback_one resetb_loopback_zero por_h porb_h porb_l mask_rev[0]
+ mask_rev[1] mask_rev[2] mask_rev[3] mask_rev[4] mask_rev[5] mask_rev[6] mask_rev[7]
+ mask_rev[8] mask_rev[9] mask_rev[10] mask_rev[11] mask_rev[12] mask_rev[13] mask_rev[14]
+ mask_rev[15] mask_rev[16] mask_rev[17] mask_rev[18] mask_rev[19] mask_rev[20] mask_rev[21]
+ mask_rev[22] mask_rev[23] mask_rev[24] mask_rev[25] mask_rev[26] mask_rev[27] mask_rev[28]
+ mask_rev[29] mask_rev[30] mask_rev[31] vssio vssd vddio vccd vert_connects_gpio_disabled_15/m2_32_14444#
+ vert_connects_gpio_disabled_27/m2_32_15194# vert_connects_gpio_disabled_27/m2_32_13800#
+ vert_connects_gpio_disabled_10/m2_32_14444# vert_connects_gpio_disabled_22/m2_32_15194#
+ vert_connects_gpio_disabled_22/m2_32_13800# vert_connects_gpio_disabled_25/m2_32_13589#
+ vert_connects_gpio_disabled_15/m2_32_15194# vert_connects_gpio_disabled_5/m2_32_14444#
+ vert_connects_gpio_disabled_15/m2_32_13800# vert_connects_gpio_disabled_20/m2_32_13589#
+ vert_connects_gpio_disabled_18/m2_32_13589# vert_connects_gpio_disabled_10/m2_32_15194#
+ vert_connects_gpio_disabled_0/m2_32_14444# vert_connects_gpio_disabled_10/m2_32_13800#
+ vert_connects_gpio_disabled_27/m2_32_14302# vert_connects_gpio_disabled_13/m2_32_13589#
+ vert_connects_gpio_disabled_22/m2_32_14302# vert_connects_gpio_disabled_26/m2_32_14673#
+ vert_connects_gpio_disabled_5/m2_32_15194# vert_connects_gpio_disabled_5/m2_32_13800#
+ vert_connects_gpio_disabled_8/m2_32_13589# vert_connects_gpio_disabled_15/m2_32_14302#
+ vert_connects_gpio_disabled_21/m2_32_14673# vert_connects_gpio_disabled_0/m2_32_15194#
+ vert_connects_gpio_disabled_0/m2_32_13800# vert_connects_gpio_disabled_19/m2_32_14673#
+ vert_connects_gpio_disabled_3/m2_32_13589# vert_connects_gpio_disabled_10/m2_32_14302#
+ vert_connects_gpio_disabled_14/m2_32_14673# vert_connects_gpio_disabled_5/m2_32_14302#
+ vert_connects_gpio_disabled_9/m2_32_14673# vert_connects_gpio_disabled_26/m2_32_14444#
+ vert_connects_gpio_disabled_0/m2_32_14302# vert_connects_gpio_disabled_4/m2_32_14673#
+ vert_connects_gpio_disabled_21/m2_32_14444# vert_connects_gpio_disabled_19/m2_32_14444#
+ vert_connects_gpio_disabled_20/m2_32_1840# vert_connects_gpio_disabled_20/m2_32_1986#
+ vert_connects_gpio_disabled_14/m2_32_14444# vert_connects_gpio_disabled_26/m2_32_15194#
+ vert_connects_gpio_disabled_26/m2_32_13800# vert_connects_gpio_disabled_21/m2_32_1840#
+ vert_connects_gpio_disabled_21/m2_32_1986# vert_connects_gpio_disabled_21/m2_32_15194#
+ vert_connects_gpio_disabled_21/m2_32_13800# vert_connects_gpio_disabled_19/m2_32_13800#
+ vert_connects_gpio_disabled_9/m2_32_14444# vert_connects_gpio_disabled_19/m2_32_15194#
+ vert_connects_gpio_disabled_22/m2_32_1840# vert_connects_gpio_disabled_24/m2_32_13589#
+ vert_connects_gpio_disabled_22/m2_32_1986# vert_connects_gpio_disabled_14/m2_32_13800#
+ vert_connects_gpio_disabled_14/m2_32_15194# vert_connects_gpio_disabled_4/m2_32_14444#
+ vert_connects_gpio_disabled_23/m2_32_1840# vert_connects_gpio_disabled_17/m2_32_13589#
+ vert_connects_gpio_disabled_23/m2_32_1986# vert_connects_gpio_disabled_26/m2_32_14302#
+ vert_connects_gpio_disabled_12/m2_32_13589# vert_connects_gpio_disabled_9/m2_32_13800#
+ vert_connects_gpio_disabled_9/m2_32_15194# vert_connects_gpio_disabled_24/m2_32_1840#
+ vert_connects_gpio_disabled_24/m2_32_1986# vert_connects_gpio_disabled_21/m2_32_14302#
+ vert_connects_gpio_disabled_19/m2_32_14302# vert_connects_gpio_disabled_25/m2_32_14673#
+ vert_connects_gpio_disabled_4/m2_32_13800# vert_connects_gpio_disabled_4/m2_32_15194#
+ vert_connects_gpio_disabled_25/m2_32_1840# vert_connects_gpio_disabled_7/m2_32_13589#
+ vert_connects_gpio_disabled_25/m2_32_1986# vert_connects_gpio_disabled_14/m2_32_14302#
+ vert_connects_gpio_disabled_20/m2_32_14673# vert_connects_gpio_disabled_18/m2_32_14673#
+ vert_connects_gpio_disabled_2/m2_32_13589# vert_connects_gpio_disabled_26/m2_32_1840#
+ vert_connects_gpio_disabled_13/m2_32_14673# vert_connects_gpio_disabled_26/m2_32_1986#
+ vert_connects_gpio_disabled_9/m2_32_14302# vert_connects_gpio_disabled_0/m2_32_1840#
+ vert_connects_gpio_disabled_0/m2_32_1986# vert_connects_gpio_disabled_27/m2_32_1840#
+ vert_connects_gpio_disabled_27/m2_32_1986# vert_connects_gpio_disabled_4/m2_32_14302#
+ vert_connects_gpio_disabled_8/m2_32_14673# vert_connects_gpio_disabled_25/m2_32_14444#
+ vert_connects_gpio_disabled_1/m2_32_1840# vert_connects_gpio_disabled_28/m2_32_1840#
+ vert_connects_gpio_disabled_1/m2_32_1986# vert_connects_gpio_disabled_28/m2_32_1986#
+ vert_connects_gpio_disabled_3/m2_32_14673# vert_connects_gpio_disabled_20/m2_32_14444#
+ gpio_drive1[15] vert_connects_gpio_disabled_20/m2_32_2132# vert_connects_gpio_disabled_18/m2_32_14444#
+ vert_connects_gpio_disabled_2/m2_32_1840# vert_connects_gpio_disabled_10/m2_32_1840#
+ vert_connects_gpio_disabled_2/m2_32_1986# vert_connects_gpio_disabled_10/m2_32_1986#
+ vert_connects_gpio_disabled_13/m2_32_14444# vert_connects_gpio_disabled_21/m2_32_2132#
+ vert_connects_gpio_disabled_25/m2_32_15194# vert_connects_gpio_disabled_3/m2_32_1840#
+ vert_connects_gpio_disabled_25/m2_32_13800# vert_connects_gpio_disabled_3/m2_32_1986#
+ vert_connects_gpio_disabled_11/m2_32_1840# vert_connects_gpio_disabled_11/m2_32_1986#
+ vert_connects_gpio_disabled_28/m2_32_13589# vert_connects_gpio_disabled_22/m2_32_2132#
+ vert_connects_gpio_disabled_20/m2_32_15194# vert_connects_gpio_disabled_20/m2_32_13800#
+ vert_connects_gpio_disabled_8/m2_32_14444# vert_connects_gpio_disabled_18/m2_32_13800#
+ vert_connects_gpio_disabled_18/m2_32_15194# vert_connects_gpio_disabled_4/m2_32_1840#
+ vert_connects_gpio_disabled_12/m2_32_1840# vert_connects_gpio_disabled_4/m2_32_1986#
+ vert_connects_gpio_disabled_23/m2_32_13589# vert_connects_gpio_disabled_12/m2_32_1986#
+ vert_connects_gpio_disabled_13/m2_32_13800# vert_connects_gpio_disabled_13/m2_32_15194#
+ vert_connects_gpio_disabled_3/m2_32_14444# vert_connects_gpio_disabled_23/m2_32_2132#
+ vert_connects_gpio_disabled_5/m2_32_1840# vert_connects_gpio_disabled_5/m2_32_1986#
+ vert_connects_gpio_disabled_13/m2_32_1840# vert_connects_gpio_disabled_16/m2_32_13589#
+ vert_connects_gpio_disabled_13/m2_32_1986# vert_connects_gpio_disabled_25/m2_32_14302#
+ vert_connects_gpio_disabled_24/m2_32_2132# vert_connects_gpio_disabled_8/m2_32_13800#
+ vert_connects_gpio_disabled_6/m2_32_1840# vert_connects_gpio_disabled_8/m2_32_15194#
+ vert_connects_gpio_disabled_11/m2_32_13589# vert_connects_gpio_disabled_14/m2_32_1840#
+ vert_connects_gpio_disabled_6/m2_32_1986# vert_connects_gpio_disabled_14/m2_32_1986#
+ vert_connects_gpio_disabled_20/m2_32_14302# vert_connects_gpio_disabled_18/m2_32_14302#
+ vert_connects_gpio_disabled_24/m2_32_14673# vert_connects_gpio_disabled_3/m2_32_15194#
+ vert_connects_gpio_disabled_25/m2_32_2132# vert_connects_gpio_disabled_3/m2_32_13800#
+ vert_connects_gpio_disabled_7/m2_32_1840# vert_connects_gpio_disabled_7/m2_32_1986#
+ vert_connects_gpio_disabled_15/m2_32_1840# vert_connects_gpio_disabled_15/m2_32_1986#
+ vert_connects_gpio_disabled_6/m2_32_13589# vert_connects_gpio_disabled_13/m2_32_14302#
+ vert_connects_gpio_disabled_17/m2_32_14673# vert_connects_gpio_disabled_26/m2_32_2132#
+ vert_connects_gpio_disabled_8/m2_32_1840# vert_connects_gpio_disabled_1/m2_32_13589#
+ vert_connects_gpio_disabled_8/m2_32_1986# vert_connects_gpio_disabled_16/m2_32_1840#
+ vert_connects_gpio_disabled_12/m2_32_14673# vert_connects_gpio_disabled_16/m2_32_1986#
+ vert_connects_gpio_disabled_8/m2_32_14302# vert_connects_gpio_disabled_0/m2_32_2132#
+ vert_connects_gpio_disabled_27/m2_32_2132# vert_connects_gpio_disabled_9/m2_32_1840#
+ vert_connects_gpio_disabled_9/m2_32_1986# vert_connects_gpio_disabled_17/m2_32_1840#
+ vert_connects_gpio_disabled_17/m2_32_1986# vert_connects_gpio_disabled_3/m2_32_14302#
+ vert_connects_gpio_disabled_7/m2_32_14673# vert_connects_gpio_disabled_1/m2_32_2132#
+ vert_connects_gpio_disabled_28/m2_32_2132# vert_connects_gpio_disabled_24/m2_32_14444#
+ vert_connects_gpio_disabled_18/m2_32_1840# vert_connects_gpio_disabled_18/m2_32_1986#
+ vert_connects_gpio_disabled_2/m2_32_14673# vert_connects_gpio_disabled_2/m2_32_2132#
+ vert_connects_gpio_disabled_10/m2_32_2132# vert_connects_gpio_disabled_17/m2_32_14444#
+ vert_connects_gpio_disabled_19/m2_32_1840# vert_connects_gpio_disabled_19/m2_32_1986#
+ vert_connects_gpio_disabled_12/m2_32_14444# vert_connects_gpio_disabled_3/m2_32_2132#
+ vert_connects_gpio_disabled_11/m2_32_2132# vert_connects_gpio_disabled_24/m2_32_15194#
+ vert_connects_gpio_disabled_24/m2_32_13800# vert_connects_gpio_disabled_27/m2_32_13589#
+ vert_connects_gpio_disabled_4/m2_32_2132# vert_connects_gpio_disabled_12/m2_32_2132#
+ vert_connects_gpio_disabled_7/m2_32_14444# vert_connects_gpio_disabled_17/m2_32_15194#
+ vert_connects_gpio_disabled_17/m2_32_13800# vert_connects_gpio_disabled_22/m2_32_13589#
+ vert_connects_gpio_disabled_5/m2_32_2132# vert_connects_gpio_disabled_2/m2_32_14444#
+ vert_connects_gpio_disabled_12/m2_32_15194# vert_connects_gpio_disabled_12/m2_32_13800#
+ vert_connects_gpio_disabled_13/m2_32_2132# vert_connects_gpio_disabled_15/m2_32_13589#
+ vert_connects_gpio_disabled_6/m2_32_2132# vert_connects_gpio_disabled_24/m2_32_14302#
+ vert_connects_gpio_disabled_14/m2_32_2132# vert_connects_gpio_disabled_28/m2_32_14673#
+ vert_connects_gpio_disabled_10/m2_32_13589# vert_connects_gpio_disabled_7/m2_32_15194#
+ vert_connects_gpio_disabled_7/m2_32_13800# vert_connects_gpio_disabled_7/m2_32_2132#
+ vert_connects_gpio_disabled_17/m2_32_14302# vert_connects_gpio_disabled_23/m2_32_14673#
+ vert_connects_gpio_disabled_2/m2_32_15194# vert_connects_gpio_disabled_15/m2_32_2132#
+ vert_connects_gpio_disabled_2/m2_32_13800# vert_connects_gpio_disabled_5/m2_32_13589#
+ vert_connects_gpio_disabled_12/m2_32_14302# vert_connects_gpio_disabled_16/m2_32_14673#
+ vert_connects_gpio_disabled_8/m2_32_2132# vert_connects_gpio_disabled_16/m2_32_2132#
+ vert_connects_gpio_disabled_0/m2_32_13589# vert_connects_gpio_disabled_11/m2_32_14673#
+ vert_connects_gpio_disabled_9/m2_32_2132# vert_connects_gpio_disabled_7/m2_32_14302#
+ vert_connects_gpio_disabled_17/m2_32_2132# vert_connects_gpio_disabled_28/m2_32_14444#
+ vert_connects_gpio_disabled_2/m2_32_14302# vert_connects_gpio_disabled_6/m2_32_14673#
+ vert_connects_gpio_disabled_18/m2_32_2132# vert_connects_gpio_disabled_23/m2_32_14444#
+ vert_connects_gpio_disabled_1/m2_32_14673# vert_connects_gpio_disabled_19/m2_32_2132#
+ vert_connects_gpio_disabled_16/m2_32_14444# vert_connects_gpio_disabled_28/m2_32_15194#
+ vert_connects_gpio_disabled_28/m2_32_13800# vert_connects_gpio_disabled_11/m2_32_14444#
+ vert_connects_gpio_disabled_23/m2_32_15194# vert_connects_gpio_disabled_23/m2_32_13800#
+ vert_connects_gpio_disabled_26/m2_32_13589# vert_connects_gpio_disabled_16/m2_32_15194#
+ vert_connects_gpio_disabled_16/m2_32_13800# vert_connects_gpio_disabled_6/m2_32_14444#
+ vert_connects_gpio_disabled_21/m2_32_13589# vert_connects_gpio_disabled_19/m2_32_13589#
+ vert_connects_gpio_disabled_11/m2_32_15194# vert_connects_gpio_disabled_11/m2_32_13800#
+ vert_connects_gpio_disabled_1/m2_32_14444# vert_connects_gpio_disabled_28/m2_32_14302#
+ vert_connects_gpio_disabled_14/m2_32_13589# vert_connects_gpio_disabled_23/m2_32_14302#
+ vert_connects_gpio_disabled_27/m2_32_14673# vert_connects_gpio_disabled_6/m2_32_15194#
+ vert_connects_gpio_disabled_6/m2_32_13800# vert_connects_gpio_disabled_9/m2_32_13589#
+ vert_connects_gpio_disabled_16/m2_32_14302# vert_connects_gpio_disabled_22/m2_32_14673#
+ vert_connects_gpio_disabled_1/m2_32_15194# vert_connects_gpio_disabled_1/m2_32_13800#
+ vert_connects_gpio_disabled_4/m2_32_13589# vert_connects_gpio_disabled_11/m2_32_14302#
+ vert_connects_gpio_disabled_15/m2_32_14673# vert_connects_gpio_disabled_10/m2_32_14673#
+ vert_connects_gpio_disabled_6/m2_32_14302# vert_connects_gpio_disabled_27/m2_32_14444#
+ vert_connects_gpio_disabled_1/m2_32_14302# vert_connects_gpio_disabled_5/m2_32_14673#
+ vert_connects_gpio_disabled_22/m2_32_14444# vert_connects_gpio_disabled_0/m2_32_14673#
Xhorz_connects_gpio_disabled_1 gpio_loopback_zero[38] gpio_pulldown[38] gpio_loopback_one[38]
+ gpio_drive0[38] gpio_drive1[38] gpio_slew[38] gpio_schmitt[38] gpio_pullup[38] gpio_out[38]
+ gpio_ie[38] gpio_oe[38] horz_connects_gpio_disabled
Xhorz_connects_gpio_disabled_2 gpio_loopback_zero[39] gpio_pulldown[39] gpio_loopback_one[39]
+ gpio_drive0[39] gpio_drive1[39] gpio_slew[39] gpio_schmitt[39] gpio_pullup[39] gpio_out[39]
+ gpio_ie[39] gpio_oe[39] horz_connects_gpio_disabled
Xhorz_connects_gpio_disabled_3 gpio_loopback_zero[40] gpio_pulldown[40] gpio_loopback_one[40]
+ gpio_drive0[40] gpio_drive1[40] gpio_slew[40] gpio_schmitt[40] gpio_pullup[40] gpio_out[40]
+ gpio_ie[40] gpio_oe[40] horz_connects_gpio_disabled
Xvert_connects_gpio_disabled_0 gpio_loopback_zero[37] gpio_drive0[37] gpio_pulldown[37]
+ gpio_schmitt[37] vert_connects_gpio_disabled_0/m2_32_14673# gpio_drive1[37] vert_connects_gpio_disabled_0/m2_32_14444#
+ vert_connects_gpio_disabled_0/m2_32_13800# vert_connects_gpio_disabled_0/m2_32_15194#
+ vert_connects_gpio_disabled_0/m2_32_14302# gpio_oe[37] gpio_out[37] vert_connects_gpio_disabled_0/m2_32_1840#
+ vert_connects_gpio_disabled_0/m2_32_1986# gpio_loopback_one[37] gpio_slew[37] vert_connects_gpio_disabled_0/m2_32_2132#
+ gpio_ie[37] vert_connects_gpio_disabled_0/m2_32_13589# gpio_pullup[37] vert_connects_gpio_disabled
Xhorz_connects_gpio_disabled_4 gpio_loopback_zero[41] gpio_pulldown[41] gpio_loopback_one[41]
+ gpio_drive0[41] gpio_drive1[41] gpio_slew[41] gpio_schmitt[41] gpio_pullup[41] gpio_out[41]
+ gpio_ie[41] gpio_oe[41] horz_connects_gpio_disabled
Xvert_connects_gpio_disabled_1 gpio_loopback_zero[36] gpio_drive0[36] gpio_pulldown[36]
+ gpio_schmitt[36] vert_connects_gpio_disabled_1/m2_32_14673# gpio_drive1[36] vert_connects_gpio_disabled_1/m2_32_14444#
+ vert_connects_gpio_disabled_1/m2_32_13800# vert_connects_gpio_disabled_1/m2_32_15194#
+ vert_connects_gpio_disabled_1/m2_32_14302# gpio_oe[36] gpio_out[36] vert_connects_gpio_disabled_1/m2_32_1840#
+ vert_connects_gpio_disabled_1/m2_32_1986# gpio_loopback_one[36] gpio_slew[36] vert_connects_gpio_disabled_1/m2_32_2132#
+ gpio_ie[36] vert_connects_gpio_disabled_1/m2_32_13589# gpio_pullup[36] vert_connects_gpio_disabled
Xhorz_connects_gpio_disabled_5 gpio_loopback_zero[42] gpio_pulldown[42] gpio_loopback_one[42]
+ gpio_drive0[42] gpio_drive1[42] gpio_slew[42] gpio_schmitt[42] gpio_pullup[42] gpio_out[42]
+ gpio_ie[42] gpio_oe[42] horz_connects_gpio_disabled
Xvert_connects_gpio_disabled_2 gpio_loopback_zero[34] gpio_drive0[34] gpio_pulldown[34]
+ gpio_schmitt[34] vert_connects_gpio_disabled_2/m2_32_14673# gpio_drive1[34] vert_connects_gpio_disabled_2/m2_32_14444#
+ vert_connects_gpio_disabled_2/m2_32_13800# vert_connects_gpio_disabled_2/m2_32_15194#
+ vert_connects_gpio_disabled_2/m2_32_14302# gpio_oe[34] gpio_out[34] vert_connects_gpio_disabled_2/m2_32_1840#
+ vert_connects_gpio_disabled_2/m2_32_1986# gpio_loopback_one[34] gpio_slew[34] vert_connects_gpio_disabled_2/m2_32_2132#
+ gpio_ie[34] vert_connects_gpio_disabled_2/m2_32_13589# gpio_pullup[34] vert_connects_gpio_disabled
Xhorz_connects_gpio_disabled_6 gpio_loopback_zero[43] gpio_pulldown[43] gpio_loopback_one[43]
+ gpio_drive0[43] gpio_drive1[43] gpio_slew[43] gpio_schmitt[43] gpio_pullup[43] gpio_out[43]
+ gpio_ie[43] gpio_oe[43] horz_connects_gpio_disabled
Xvert_connects_gpio_disabled_3 gpio_loopback_zero[33] gpio_drive0[33] gpio_pulldown[33]
+ gpio_schmitt[33] vert_connects_gpio_disabled_3/m2_32_14673# gpio_drive1[33] vert_connects_gpio_disabled_3/m2_32_14444#
+ vert_connects_gpio_disabled_3/m2_32_13800# vert_connects_gpio_disabled_3/m2_32_15194#
+ vert_connects_gpio_disabled_3/m2_32_14302# gpio_oe[33] gpio_out[33] vert_connects_gpio_disabled_3/m2_32_1840#
+ vert_connects_gpio_disabled_3/m2_32_1986# gpio_loopback_one[33] gpio_slew[33] vert_connects_gpio_disabled_3/m2_32_2132#
+ gpio_ie[33] vert_connects_gpio_disabled_3/m2_32_13589# gpio_pullup[33] vert_connects_gpio_disabled
Xvert_connects_gpio_disabled_20 gpio_loopback_zero[7] gpio_drive0[7] gpio_pulldown[7]
+ gpio_schmitt[7] vert_connects_gpio_disabled_20/m2_32_14673# gpio_drive1[7] vert_connects_gpio_disabled_20/m2_32_14444#
+ vert_connects_gpio_disabled_20/m2_32_13800# vert_connects_gpio_disabled_20/m2_32_15194#
+ vert_connects_gpio_disabled_20/m2_32_14302# gpio_oe[7] gpio_out[7] vert_connects_gpio_disabled_20/m2_32_1840#
+ vert_connects_gpio_disabled_20/m2_32_1986# gpio_loopback_one[7] gpio_slew[7] vert_connects_gpio_disabled_20/m2_32_2132#
+ gpio_ie[7] vert_connects_gpio_disabled_20/m2_32_13589# gpio_pullup[7] vert_connects_gpio_disabled
Xhorz_connects_gpio_disabled_7 gpio_loopback_zero[15] gpio_pulldown[15] gpio_loopback_one[15]
+ gpio_drive0[15] gpio_drive1[15] gpio_slew[15] gpio_schmitt[15] gpio_pullup[15] gpio_out[15]
+ gpio_ie[15] gpio_oe[15] horz_connects_gpio_disabled
Xvert_connects_gpio_disabled_4 gpio_loopback_zero[32] gpio_drive0[32] gpio_pulldown[32]
+ gpio_schmitt[32] vert_connects_gpio_disabled_4/m2_32_14673# gpio_drive1[32] vert_connects_gpio_disabled_4/m2_32_14444#
+ vert_connects_gpio_disabled_4/m2_32_13800# vert_connects_gpio_disabled_4/m2_32_15194#
+ vert_connects_gpio_disabled_4/m2_32_14302# gpio_oe[32] gpio_out[32] vert_connects_gpio_disabled_4/m2_32_1840#
+ vert_connects_gpio_disabled_4/m2_32_1986# gpio_loopback_one[32] gpio_slew[32] vert_connects_gpio_disabled_4/m2_32_2132#
+ gpio_ie[32] vert_connects_gpio_disabled_4/m2_32_13589# gpio_pullup[32] vert_connects_gpio_disabled
Xvert_connects_gpio_disabled_10 gpio_loopback_zero[26] gpio_drive0[26] gpio_pulldown[26]
+ gpio_schmitt[26] vert_connects_gpio_disabled_10/m2_32_14673# gpio_drive1[26] vert_connects_gpio_disabled_10/m2_32_14444#
+ vert_connects_gpio_disabled_10/m2_32_13800# vert_connects_gpio_disabled_10/m2_32_15194#
+ vert_connects_gpio_disabled_10/m2_32_14302# gpio_oe[26] gpio_out[26] vert_connects_gpio_disabled_10/m2_32_1840#
+ vert_connects_gpio_disabled_10/m2_32_1986# gpio_loopback_one[26] gpio_slew[26] vert_connects_gpio_disabled_10/m2_32_2132#
+ gpio_ie[26] vert_connects_gpio_disabled_10/m2_32_13589# gpio_pullup[26] vert_connects_gpio_disabled
Xvert_connects_gpio_disabled_21 gpio_loopback_zero[8] gpio_drive0[8] gpio_pulldown[8]
+ gpio_schmitt[8] vert_connects_gpio_disabled_21/m2_32_14673# gpio_drive1[8] vert_connects_gpio_disabled_21/m2_32_14444#
+ vert_connects_gpio_disabled_21/m2_32_13800# vert_connects_gpio_disabled_21/m2_32_15194#
+ vert_connects_gpio_disabled_21/m2_32_14302# gpio_oe[8] gpio_out[8] vert_connects_gpio_disabled_21/m2_32_1840#
+ vert_connects_gpio_disabled_21/m2_32_1986# gpio_loopback_one[8] gpio_slew[8] vert_connects_gpio_disabled_21/m2_32_2132#
+ gpio_ie[8] vert_connects_gpio_disabled_21/m2_32_13589# gpio_pullup[8] vert_connects_gpio_disabled
Xhorz_connects_gpio_disabled_8 gpio_loopback_zero[16] gpio_pulldown[16] gpio_loopback_one[16]
+ gpio_drive0[16] gpio_drive1[16] gpio_slew[16] gpio_schmitt[16] gpio_pullup[16] gpio_out[16]
+ gpio_ie[16] gpio_oe[16] horz_connects_gpio_disabled
Xhorz_connects_gpio_disabled_9 gpio_loopback_zero[17] gpio_pulldown[17] gpio_loopback_one[17]
+ gpio_drive0[17] gpio_drive1[17] gpio_slew[17] gpio_schmitt[17] gpio_pullup[17] gpio_out[17]
+ gpio_ie[17] gpio_oe[17] horz_connects_gpio_disabled
Xhorz_connects_gpio_disabled_10 gpio_loopback_zero[18] gpio_pulldown[18] gpio_loopback_one[18]
+ gpio_drive0[18] gpio_drive1[18] gpio_slew[18] gpio_schmitt[18] gpio_pullup[18] gpio_out[18]
+ gpio_ie[18] gpio_oe[18] horz_connects_gpio_disabled
Xvert_connects_gpio_disabled_5 gpio_loopback_zero[31] gpio_drive0[31] gpio_pulldown[31]
+ gpio_schmitt[31] vert_connects_gpio_disabled_5/m2_32_14673# gpio_drive1[31] vert_connects_gpio_disabled_5/m2_32_14444#
+ vert_connects_gpio_disabled_5/m2_32_13800# vert_connects_gpio_disabled_5/m2_32_15194#
+ vert_connects_gpio_disabled_5/m2_32_14302# gpio_oe[31] gpio_out[31] vert_connects_gpio_disabled_5/m2_32_1840#
+ vert_connects_gpio_disabled_5/m2_32_1986# gpio_loopback_one[31] gpio_slew[31] vert_connects_gpio_disabled_5/m2_32_2132#
+ gpio_ie[31] vert_connects_gpio_disabled_5/m2_32_13589# gpio_pullup[31] vert_connects_gpio_disabled
Xvert_connects_gpio_disabled_11 gpio_loopback_zero[25] gpio_drive0[25] gpio_pulldown[25]
+ gpio_schmitt[25] vert_connects_gpio_disabled_11/m2_32_14673# gpio_drive1[25] vert_connects_gpio_disabled_11/m2_32_14444#
+ vert_connects_gpio_disabled_11/m2_32_13800# vert_connects_gpio_disabled_11/m2_32_15194#
+ vert_connects_gpio_disabled_11/m2_32_14302# gpio_oe[25] gpio_out[25] vert_connects_gpio_disabled_11/m2_32_1840#
+ vert_connects_gpio_disabled_11/m2_32_1986# gpio_loopback_one[25] gpio_slew[25] vert_connects_gpio_disabled_11/m2_32_2132#
+ gpio_ie[25] vert_connects_gpio_disabled_11/m2_32_13589# gpio_pullup[25] vert_connects_gpio_disabled
Xvert_connects_gpio_disabled_22 gpio_loopback_zero[9] gpio_drive0[9] gpio_pulldown[9]
+ gpio_schmitt[9] vert_connects_gpio_disabled_22/m2_32_14673# gpio_drive1[9] vert_connects_gpio_disabled_22/m2_32_14444#
+ vert_connects_gpio_disabled_22/m2_32_13800# vert_connects_gpio_disabled_22/m2_32_15194#
+ vert_connects_gpio_disabled_22/m2_32_14302# gpio_oe[9] gpio_out[9] vert_connects_gpio_disabled_22/m2_32_1840#
+ vert_connects_gpio_disabled_22/m2_32_1986# gpio_loopback_one[9] gpio_slew[9] vert_connects_gpio_disabled_22/m2_32_2132#
+ gpio_ie[9] vert_connects_gpio_disabled_22/m2_32_13589# gpio_pullup[9] vert_connects_gpio_disabled
Xhorz_connects_gpio_disabled_11 gpio_loopback_zero[19] gpio_pulldown[19] gpio_loopback_one[19]
+ gpio_drive0[19] gpio_drive1[19] gpio_slew[19] gpio_schmitt[19] gpio_pullup[19] gpio_out[19]
+ gpio_ie[19] gpio_oe[19] horz_connects_gpio_disabled
Xvert_connects_gpio_disabled_6 gpio_loopback_zero[30] gpio_drive0[30] gpio_pulldown[30]
+ gpio_schmitt[30] vert_connects_gpio_disabled_6/m2_32_14673# gpio_drive1[30] vert_connects_gpio_disabled_6/m2_32_14444#
+ vert_connects_gpio_disabled_6/m2_32_13800# vert_connects_gpio_disabled_6/m2_32_15194#
+ vert_connects_gpio_disabled_6/m2_32_14302# gpio_oe[30] gpio_out[30] vert_connects_gpio_disabled_6/m2_32_1840#
+ vert_connects_gpio_disabled_6/m2_32_1986# gpio_loopback_one[30] gpio_slew[30] vert_connects_gpio_disabled_6/m2_32_2132#
+ gpio_ie[30] vert_connects_gpio_disabled_6/m2_32_13589# gpio_pullup[30] vert_connects_gpio_disabled
Xvert_connects_gpio_disabled_7 gpio_loopback_zero[29] gpio_drive0[29] gpio_pulldown[29]
+ gpio_schmitt[29] vert_connects_gpio_disabled_7/m2_32_14673# gpio_drive1[29] vert_connects_gpio_disabled_7/m2_32_14444#
+ vert_connects_gpio_disabled_7/m2_32_13800# vert_connects_gpio_disabled_7/m2_32_15194#
+ vert_connects_gpio_disabled_7/m2_32_14302# gpio_oe[29] gpio_out[29] vert_connects_gpio_disabled_7/m2_32_1840#
+ vert_connects_gpio_disabled_7/m2_32_1986# gpio_loopback_one[29] gpio_slew[29] vert_connects_gpio_disabled_7/m2_32_2132#
+ gpio_ie[29] vert_connects_gpio_disabled_7/m2_32_13589# gpio_pullup[29] vert_connects_gpio_disabled
Xvert_connects_gpio_disabled_12 gpio_loopback_zero[24] gpio_drive0[24] gpio_pulldown[24]
+ gpio_schmitt[24] vert_connects_gpio_disabled_12/m2_32_14673# gpio_drive1[24] vert_connects_gpio_disabled_12/m2_32_14444#
+ vert_connects_gpio_disabled_12/m2_32_13800# vert_connects_gpio_disabled_12/m2_32_15194#
+ vert_connects_gpio_disabled_12/m2_32_14302# gpio_oe[24] gpio_out[24] vert_connects_gpio_disabled_12/m2_32_1840#
+ vert_connects_gpio_disabled_12/m2_32_1986# gpio_loopback_one[24] gpio_slew[24] vert_connects_gpio_disabled_12/m2_32_2132#
+ gpio_ie[24] vert_connects_gpio_disabled_12/m2_32_13589# gpio_pullup[24] vert_connects_gpio_disabled
Xvert_connects_gpio_disabled_23 gpio_loopback_zero[10] gpio_drive0[10] gpio_pulldown[10]
+ gpio_schmitt[10] vert_connects_gpio_disabled_23/m2_32_14673# gpio_drive1[10] vert_connects_gpio_disabled_23/m2_32_14444#
+ vert_connects_gpio_disabled_23/m2_32_13800# vert_connects_gpio_disabled_23/m2_32_15194#
+ vert_connects_gpio_disabled_23/m2_32_14302# gpio_oe[10] gpio_out[10] vert_connects_gpio_disabled_23/m2_32_1840#
+ vert_connects_gpio_disabled_23/m2_32_1986# gpio_loopback_one[10] gpio_slew[10] vert_connects_gpio_disabled_23/m2_32_2132#
+ gpio_ie[10] vert_connects_gpio_disabled_23/m2_32_13589# gpio_pullup[10] vert_connects_gpio_disabled
Xhorz_connects_gpio_disabled_12 gpio_loopback_zero[20] gpio_pulldown[20] gpio_loopback_one[20]
+ gpio_drive0[20] gpio_drive1[20] gpio_slew[20] gpio_schmitt[20] gpio_pullup[20] gpio_out[20]
+ gpio_ie[20] gpio_oe[20] horz_connects_gpio_disabled
Xhorz_connects_gpio_disabled_13 gpio_loopback_zero[21] gpio_pulldown[21] gpio_loopback_one[21]
+ gpio_drive0[21] gpio_drive1[21] gpio_slew[21] gpio_schmitt[21] gpio_pullup[21] gpio_out[21]
+ gpio_ie[21] gpio_oe[21] horz_connects_gpio_disabled
Xvert_connects_gpio_disabled_8 gpio_loopback_zero[28] gpio_drive0[28] gpio_pulldown[28]
+ gpio_schmitt[28] vert_connects_gpio_disabled_8/m2_32_14673# gpio_drive1[28] vert_connects_gpio_disabled_8/m2_32_14444#
+ vert_connects_gpio_disabled_8/m2_32_13800# vert_connects_gpio_disabled_8/m2_32_15194#
+ vert_connects_gpio_disabled_8/m2_32_14302# gpio_oe[28] gpio_out[28] vert_connects_gpio_disabled_8/m2_32_1840#
+ vert_connects_gpio_disabled_8/m2_32_1986# gpio_loopback_one[28] gpio_slew[28] vert_connects_gpio_disabled_8/m2_32_2132#
+ gpio_ie[28] vert_connects_gpio_disabled_8/m2_32_13589# gpio_pullup[28] vert_connects_gpio_disabled
Xvert_connects_gpio_disabled_13 gpio_loopback_zero[0] gpio_drive0[0] gpio_pulldown[0]
+ gpio_schmitt[0] vert_connects_gpio_disabled_13/m2_32_14673# gpio_drive1[0] vert_connects_gpio_disabled_13/m2_32_14444#
+ vert_connects_gpio_disabled_13/m2_32_13800# vert_connects_gpio_disabled_13/m2_32_15194#
+ vert_connects_gpio_disabled_13/m2_32_14302# gpio_oe[0] gpio_out[0] vert_connects_gpio_disabled_13/m2_32_1840#
+ vert_connects_gpio_disabled_13/m2_32_1986# gpio_loopback_one[0] gpio_slew[0] vert_connects_gpio_disabled_13/m2_32_2132#
+ gpio_ie[0] vert_connects_gpio_disabled_13/m2_32_13589# gpio_pullup[0] vert_connects_gpio_disabled
Xvert_connects_gpio_disabled_24 gpio_loopback_zero[11] gpio_drive0[11] gpio_pulldown[11]
+ gpio_schmitt[11] vert_connects_gpio_disabled_24/m2_32_14673# gpio_drive1[11] vert_connects_gpio_disabled_24/m2_32_14444#
+ vert_connects_gpio_disabled_24/m2_32_13800# vert_connects_gpio_disabled_24/m2_32_15194#
+ vert_connects_gpio_disabled_24/m2_32_14302# gpio_oe[11] gpio_out[11] vert_connects_gpio_disabled_24/m2_32_1840#
+ vert_connects_gpio_disabled_24/m2_32_1986# gpio_loopback_one[11] gpio_slew[11] vert_connects_gpio_disabled_24/m2_32_2132#
+ gpio_ie[11] vert_connects_gpio_disabled_24/m2_32_13589# gpio_pullup[11] vert_connects_gpio_disabled
Xhorz_connects_gpio_disabled_14 gpio_loopback_zero[22] gpio_pulldown[22] gpio_loopback_one[22]
+ gpio_drive0[22] gpio_drive1[22] gpio_slew[22] gpio_schmitt[22] gpio_pullup[22] gpio_out[22]
+ gpio_ie[22] gpio_oe[22] horz_connects_gpio_disabled
Xvert_connects_gpio_disabled_9 gpio_loopback_zero[27] gpio_drive0[27] gpio_pulldown[27]
+ gpio_schmitt[27] vert_connects_gpio_disabled_9/m2_32_14673# gpio_drive1[27] vert_connects_gpio_disabled_9/m2_32_14444#
+ vert_connects_gpio_disabled_9/m2_32_13800# vert_connects_gpio_disabled_9/m2_32_15194#
+ vert_connects_gpio_disabled_9/m2_32_14302# gpio_oe[27] gpio_out[27] vert_connects_gpio_disabled_9/m2_32_1840#
+ vert_connects_gpio_disabled_9/m2_32_1986# gpio_loopback_one[27] gpio_slew[27] vert_connects_gpio_disabled_9/m2_32_2132#
+ gpio_ie[27] vert_connects_gpio_disabled_9/m2_32_13589# gpio_pullup[27] vert_connects_gpio_disabled
Xvert_connects_gpio_disabled_14 gpio_loopback_zero[1] gpio_drive0[1] gpio_pulldown[1]
+ gpio_schmitt[1] vert_connects_gpio_disabled_14/m2_32_14673# gpio_drive1[1] vert_connects_gpio_disabled_14/m2_32_14444#
+ vert_connects_gpio_disabled_14/m2_32_13800# vert_connects_gpio_disabled_14/m2_32_15194#
+ vert_connects_gpio_disabled_14/m2_32_14302# gpio_oe[1] gpio_out[1] vert_connects_gpio_disabled_14/m2_32_1840#
+ vert_connects_gpio_disabled_14/m2_32_1986# gpio_loopback_one[1] gpio_slew[1] vert_connects_gpio_disabled_14/m2_32_2132#
+ gpio_ie[1] vert_connects_gpio_disabled_14/m2_32_13589# gpio_pullup[1] vert_connects_gpio_disabled
Xvert_connects_gpio_disabled_25 gpio_loopback_zero[12] gpio_drive0[12] gpio_pulldown[12]
+ gpio_schmitt[12] vert_connects_gpio_disabled_25/m2_32_14673# gpio_drive1[12] vert_connects_gpio_disabled_25/m2_32_14444#
+ vert_connects_gpio_disabled_25/m2_32_13800# vert_connects_gpio_disabled_25/m2_32_15194#
+ vert_connects_gpio_disabled_25/m2_32_14302# gpio_oe[12] gpio_out[12] vert_connects_gpio_disabled_25/m2_32_1840#
+ vert_connects_gpio_disabled_25/m2_32_1986# gpio_loopback_one[12] gpio_slew[12] vert_connects_gpio_disabled_25/m2_32_2132#
+ gpio_ie[12] vert_connects_gpio_disabled_25/m2_32_13589# gpio_pullup[12] vert_connects_gpio_disabled
Xhorz_connects_gpio_disabled_15 gpio_loopback_zero[23] gpio_pulldown[23] gpio_loopback_one[23]
+ gpio_drive0[23] gpio_drive1[23] gpio_slew[23] gpio_schmitt[23] gpio_pullup[23] gpio_out[23]
+ gpio_ie[23] gpio_oe[23] horz_connects_gpio_disabled
Xvert_connects_gpio_disabled_15 gpio_loopback_zero[2] gpio_drive0[2] gpio_pulldown[2]
+ gpio_schmitt[2] vert_connects_gpio_disabled_15/m2_32_14673# gpio_drive1[2] vert_connects_gpio_disabled_15/m2_32_14444#
+ vert_connects_gpio_disabled_15/m2_32_13800# vert_connects_gpio_disabled_15/m2_32_15194#
+ vert_connects_gpio_disabled_15/m2_32_14302# gpio_oe[2] gpio_out[2] vert_connects_gpio_disabled_15/m2_32_1840#
+ vert_connects_gpio_disabled_15/m2_32_1986# gpio_loopback_one[2] gpio_slew[2] vert_connects_gpio_disabled_15/m2_32_2132#
+ gpio_ie[2] vert_connects_gpio_disabled_15/m2_32_13589# gpio_pullup[2] vert_connects_gpio_disabled
Xvert_connects_gpio_disabled_26 gpio_loopback_zero[13] gpio_drive0[13] gpio_pulldown[13]
+ gpio_schmitt[13] vert_connects_gpio_disabled_26/m2_32_14673# gpio_drive1[13] vert_connects_gpio_disabled_26/m2_32_14444#
+ vert_connects_gpio_disabled_26/m2_32_13800# vert_connects_gpio_disabled_26/m2_32_15194#
+ vert_connects_gpio_disabled_26/m2_32_14302# gpio_oe[13] gpio_out[13] vert_connects_gpio_disabled_26/m2_32_1840#
+ vert_connects_gpio_disabled_26/m2_32_1986# gpio_loopback_one[13] gpio_slew[13] vert_connects_gpio_disabled_26/m2_32_2132#
+ gpio_ie[13] vert_connects_gpio_disabled_26/m2_32_13589# gpio_pullup[13] vert_connects_gpio_disabled
Xvert_connects_gpio_disabled_16 gpio_loopback_zero[3] gpio_drive0[3] gpio_pulldown[3]
+ gpio_schmitt[3] vert_connects_gpio_disabled_16/m2_32_14673# gpio_drive1[3] vert_connects_gpio_disabled_16/m2_32_14444#
+ vert_connects_gpio_disabled_16/m2_32_13800# vert_connects_gpio_disabled_16/m2_32_15194#
+ vert_connects_gpio_disabled_16/m2_32_14302# gpio_oe[3] gpio_out[3] vert_connects_gpio_disabled_16/m2_32_1840#
+ vert_connects_gpio_disabled_16/m2_32_1986# gpio_loopback_one[3] gpio_slew[3] vert_connects_gpio_disabled_16/m2_32_2132#
+ gpio_ie[3] vert_connects_gpio_disabled_16/m2_32_13589# gpio_pullup[3] vert_connects_gpio_disabled
Xvert_connects_gpio_disabled_27 gpio_loopback_zero[14] gpio_drive0[14] gpio_pulldown[14]
+ gpio_schmitt[14] vert_connects_gpio_disabled_27/m2_32_14673# gpio_drive1[14] vert_connects_gpio_disabled_27/m2_32_14444#
+ vert_connects_gpio_disabled_27/m2_32_13800# vert_connects_gpio_disabled_27/m2_32_15194#
+ vert_connects_gpio_disabled_27/m2_32_14302# gpio_oe[14] gpio_out[14] vert_connects_gpio_disabled_27/m2_32_1840#
+ vert_connects_gpio_disabled_27/m2_32_1986# gpio_loopback_one[14] gpio_slew[14] vert_connects_gpio_disabled_27/m2_32_2132#
+ gpio_ie[14] vert_connects_gpio_disabled_27/m2_32_13589# gpio_pullup[14] vert_connects_gpio_disabled
Xvert_connects_gpio_disabled_17 gpio_loopback_zero[4] gpio_drive0[4] gpio_pulldown[4]
+ gpio_schmitt[4] vert_connects_gpio_disabled_17/m2_32_14673# gpio_drive1[4] vert_connects_gpio_disabled_17/m2_32_14444#
+ vert_connects_gpio_disabled_17/m2_32_13800# vert_connects_gpio_disabled_17/m2_32_15194#
+ vert_connects_gpio_disabled_17/m2_32_14302# gpio_oe[4] gpio_out[4] vert_connects_gpio_disabled_17/m2_32_1840#
+ vert_connects_gpio_disabled_17/m2_32_1986# gpio_loopback_one[4] gpio_slew[4] vert_connects_gpio_disabled_17/m2_32_2132#
+ gpio_ie[4] vert_connects_gpio_disabled_17/m2_32_13589# gpio_pullup[4] vert_connects_gpio_disabled
Xvert_connects_gpio_disabled_18 gpio_loopback_zero[5] gpio_drive0[5] gpio_pulldown[5]
+ gpio_schmitt[5] vert_connects_gpio_disabled_18/m2_32_14673# gpio_drive1[5] vert_connects_gpio_disabled_18/m2_32_14444#
+ vert_connects_gpio_disabled_18/m2_32_13800# vert_connects_gpio_disabled_18/m2_32_15194#
+ vert_connects_gpio_disabled_18/m2_32_14302# gpio_oe[5] gpio_out[5] vert_connects_gpio_disabled_18/m2_32_1840#
+ vert_connects_gpio_disabled_18/m2_32_1986# gpio_loopback_one[5] gpio_slew[5] vert_connects_gpio_disabled_18/m2_32_2132#
+ gpio_ie[5] vert_connects_gpio_disabled_18/m2_32_13589# gpio_pullup[5] vert_connects_gpio_disabled
Xvert_connects_gpio_disabled_28 gpio_loopback_zero[35] gpio_drive0[35] gpio_pulldown[35]
+ gpio_schmitt[35] vert_connects_gpio_disabled_28/m2_32_14673# gpio_drive1[35] vert_connects_gpio_disabled_28/m2_32_14444#
+ vert_connects_gpio_disabled_28/m2_32_13800# vert_connects_gpio_disabled_28/m2_32_15194#
+ vert_connects_gpio_disabled_28/m2_32_14302# gpio_oe[35] gpio_out[35] vert_connects_gpio_disabled_28/m2_32_1840#
+ vert_connects_gpio_disabled_28/m2_32_1986# gpio_loopback_one[35] gpio_slew[35] vert_connects_gpio_disabled_28/m2_32_2132#
+ gpio_ie[35] vert_connects_gpio_disabled_28/m2_32_13589# gpio_pullup[35] vert_connects_gpio_disabled
Xvert_connects_gpio_disabled_19 gpio_loopback_zero[6] gpio_drive0[6] gpio_pulldown[6]
+ gpio_schmitt[6] vert_connects_gpio_disabled_19/m2_32_14673# gpio_drive1[6] vert_connects_gpio_disabled_19/m2_32_14444#
+ vert_connects_gpio_disabled_19/m2_32_13800# vert_connects_gpio_disabled_19/m2_32_15194#
+ vert_connects_gpio_disabled_19/m2_32_14302# gpio_oe[6] gpio_out[6] vert_connects_gpio_disabled_19/m2_32_1840#
+ vert_connects_gpio_disabled_19/m2_32_1986# gpio_loopback_one[6] gpio_slew[6] vert_connects_gpio_disabled_19/m2_32_2132#
+ gpio_ie[6] vert_connects_gpio_disabled_19/m2_32_13589# gpio_pullup[6] vert_connects_gpio_disabled
R0 resetb_pulldown resetb_loopback_zero 0.000000
R1 resetb_pullup resetb_loopback_one 0.000000
.ends

.subckt openframe_project_wrapper gpio_in[38] gpio_in[40] gpio_oe[40] gpio_in[39]
+ gpio_oe[39] gpio_in[41] gpio_out[41] gpio_ie[41] gpio_oe[41] gpio_in[42] gpio_out[42]
+ gpio_ie[42] gpio_oe[42] gpio_drive0[38] gpio_drive1[38] gpio_in[43] gpio_ie[38]
+ gpio_out[38] gpio_oe[38] gpio_pulldown[38] gpio_pullup[38] gpio_schmitt[38] gpio_slew[38]
+ gpio_schmitt[42] gpio_pullup[42] gpio_drive0[42] gpio_drive1[42] gpio_pulldown[42]
+ gpio_slew[42] gpio_schmitt[41] gpio_pullup[41] gpio_drive0[41] gpio_drive1[41] gpio_pulldown[41]
+ gpio_slew[41] gpio_schmitt[40] gpio_pullup[40] gpio_drive0[40] gpio_drive1[40] gpio_pulldown[40]
+ gpio_ie[40] gpio_slew[40] gpio_out[40] gpio_schmitt[39] gpio_pullup[39] gpio_drive0[39]
+ gpio_drive1[39] gpio_pulldown[39] gpio_ie[39] gpio_slew[39] gpio_out[39] gpio_out[43]
+ gpio_slew[43] gpio_ie[43] gpio_pulldown[43] gpio_drive1[43] gpio_drive0[43] gpio_pullup[43]
+ gpio_schmitt[43] gpio_oe[43] gpio_drive0[30] gpio_drive0[0] gpio_drive0[5] gpio_drive1[5]
+ gpio_drive0[6] gpio_drive1[6] gpio_drive0[7] gpio_drive1[7] gpio_drive0[8] gpio_drive1[8]
+ gpio_drive0[9] gpio_drive1[9] gpio_drive1[0] gpio_drive0[10] gpio_drive1[10] gpio_drive0[11]
+ gpio_drive1[11] gpio_drive0[12] gpio_drive1[12] gpio_drive0[13] gpio_drive1[13]
+ gpio_drive0[14] gpio_drive1[14] gpio_drive0[1] gpio_drive0[15] gpio_drive1[15] gpio_drive0[16]
+ gpio_drive1[16] gpio_drive0[17] gpio_drive1[17] gpio_drive0[18] gpio_drive1[18]
+ gpio_drive0[19] gpio_drive1[1] gpio_drive0[20] gpio_drive1[20] gpio_drive0[21] gpio_drive1[21]
+ gpio_drive0[22] gpio_drive1[22] gpio_drive0[23] gpio_drive1[23] gpio_drive0[24]
+ gpio_drive1[24] gpio_drive0[2] gpio_drive1[25] gpio_drive0[25] gpio_drive0[26] gpio_drive1[26]
+ gpio_drive0[27] gpio_drive1[27] gpio_drive0[28] gpio_drive1[28] gpio_drive0[29]
+ gpio_drive1[29] gpio_drive1[2] gpio_drive1[30] gpio_drive0[31] gpio_drive1[31] gpio_drive0[32]
+ gpio_drive1[32] gpio_drive0[33] gpio_drive1[33] gpio_drive0[34] gpio_drive1[34]
+ gpio_drive0[3] gpio_drive0[35] gpio_drive1[35] gpio_drive0[36] gpio_drive1[36] gpio_drive0[37]
+ gpio_drive1[37] gpio_drive1[3] gpio_drive0[4] gpio_drive1[4] gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[34] gpio_in[35] gpio_in[36]
+ gpio_in[37] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_ie[0] gpio_ie[10] gpio_ie[11] gpio_ie[12] gpio_ie[13] gpio_ie[14] gpio_ie[15]
+ gpio_ie[16] gpio_ie[17] gpio_ie[18] gpio_ie[19] gpio_ie[1] gpio_ie[20] gpio_ie[21]
+ gpio_ie[22] gpio_ie[23] gpio_ie[24] gpio_ie[25] gpio_ie[26] gpio_ie[27] gpio_ie[28]
+ gpio_ie[29] gpio_ie[2] gpio_ie[30] gpio_ie[31] gpio_ie[32] gpio_ie[33] gpio_ie[34]
+ gpio_ie[35] gpio_ie[36] gpio_ie[37] gpio_ie[3] gpio_ie[4] gpio_ie[5] gpio_ie[6]
+ gpio_ie[7] gpio_ie[8] gpio_ie[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[34] gpio_out[35] gpio_out[36] gpio_out[37] gpio_out[3]
+ gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] gpio_oe[0]
+ gpio_oe[10] gpio_oe[11] gpio_oe[12] gpio_oe[13] gpio_oe[14] gpio_oe[15] gpio_oe[16]
+ gpio_oe[17] gpio_oe[18] gpio_oe[19] gpio_oe[1] gpio_oe[20] gpio_oe[21] gpio_oe[22]
+ gpio_oe[23] gpio_oe[24] gpio_oe[25] gpio_oe[26] gpio_oe[27] gpio_oe[28] gpio_oe[29]
+ gpio_oe[2] gpio_oe[30] gpio_oe[31] gpio_oe[32] gpio_oe[33] gpio_oe[34] gpio_oe[35]
+ gpio_oe[36] gpio_oe[37] gpio_oe[3] gpio_oe[4] gpio_oe[5] gpio_oe[6] gpio_oe[7] gpio_oe[8]
+ gpio_oe[9] gpio_pulldown[0] gpio_pulldown[10] gpio_pulldown[11] gpio_pulldown[12]
+ gpio_pulldown[13] gpio_pulldown[14] gpio_pulldown[15] gpio_pulldown[16] gpio_pulldown[17]
+ gpio_pulldown[18] gpio_pulldown[19] gpio_pulldown[1] gpio_pulldown[20] gpio_pulldown[21]
+ gpio_pulldown[22] gpio_pulldown[23] gpio_pulldown[24] gpio_pulldown[25] gpio_pulldown[26]
+ gpio_pulldown[27] gpio_pulldown[28] gpio_pulldown[29] gpio_pulldown[2] gpio_pulldown[30]
+ gpio_pulldown[31] gpio_pulldown[32] gpio_pulldown[33] gpio_pulldown[34] gpio_pulldown[35]
+ gpio_pulldown[36] gpio_pulldown[37] gpio_pulldown[3] gpio_pulldown[4] gpio_pulldown[5]
+ gpio_pulldown[6] gpio_pulldown[7] gpio_pulldown[8] gpio_pulldown[9] gpio_pullup[0]
+ gpio_pullup[10] gpio_pullup[11] gpio_pullup[12] gpio_pullup[13] gpio_pullup[14]
+ gpio_pullup[15] gpio_pullup[16] gpio_pullup[17] gpio_pullup[18] gpio_pullup[19]
+ gpio_pullup[1] gpio_pullup[20] gpio_pullup[21] gpio_pullup[22] gpio_pullup[23] gpio_pullup[24]
+ gpio_pullup[25] gpio_pullup[26] gpio_pullup[27] gpio_pullup[28] gpio_pullup[29]
+ gpio_pullup[2] gpio_pullup[30] gpio_pullup[31] gpio_pullup[32] gpio_pullup[33] gpio_pullup[34]
+ gpio_pullup[35] gpio_pullup[36] gpio_pullup[37] gpio_pullup[3] gpio_pullup[4] gpio_pullup[5]
+ gpio_pullup[6] gpio_pullup[7] gpio_pullup[8] gpio_pullup[9] gpio_schmitt[0] gpio_schmitt[10]
+ gpio_schmitt[11] gpio_schmitt[12] gpio_schmitt[13] gpio_schmitt[14] gpio_schmitt[15]
+ gpio_schmitt[16] gpio_schmitt[17] gpio_schmitt[18] gpio_schmitt[19] gpio_schmitt[1]
+ gpio_schmitt[20] gpio_schmitt[21] gpio_schmitt[22] gpio_schmitt[23] gpio_schmitt[24]
+ gpio_schmitt[25] gpio_schmitt[26] gpio_schmitt[27] gpio_schmitt[28] gpio_schmitt[29]
+ gpio_schmitt[2] gpio_schmitt[30] gpio_schmitt[31] gpio_schmitt[32] gpio_schmitt[33]
+ gpio_schmitt[34] gpio_schmitt[35] gpio_schmitt[36] gpio_schmitt[37] gpio_schmitt[3]
+ gpio_schmitt[4] gpio_schmitt[5] gpio_schmitt[6] gpio_schmitt[7] gpio_schmitt[8]
+ gpio_schmitt[9] gpio_slew[0] gpio_slew[10] gpio_slew[11] gpio_slew[12] gpio_slew[13]
+ gpio_slew[14] gpio_slew[15] gpio_slew[16] gpio_slew[17] gpio_slew[18] gpio_slew[19]
+ gpio_slew[1] gpio_slew[20] gpio_slew[21] gpio_slew[22] gpio_slew[23] gpio_slew[24]
+ gpio_slew[25] gpio_slew[26] gpio_slew[27] gpio_slew[28] gpio_slew[29] gpio_slew[2]
+ gpio_slew[30] gpio_slew[31] gpio_slew[32] gpio_slew[33] gpio_slew[34] gpio_slew[35]
+ gpio_slew[36] gpio_slew[37] gpio_slew[3] gpio_slew[4] gpio_slew[5] gpio_slew[6]
+ gpio_slew[7] gpio_slew[8] gpio_slew[9] resetb_core gpio_ana[0] gpio_ana[1] gpio_ana[2]
+ gpio_ana[3] gpio_ana[4] gpio_ana[5] gpio_ana[6] gpio_ana[7] gpio_ana[8] gpio_ana[9]
+ gpio_ana[10] gpio_ana[11] gpio_ana[12] gpio_ana[13] gpio_ana[14] gpio_ana[15] gpio_ana[16]
+ gpio_ana[17] gpio_ana[18] gpio_ana[19] gpio_ana[20] gpio_ana[21] gpio_ana[22] gpio_ana[23]
+ gpio_ana[24] gpio_ana[25] gpio_ana[26] gpio_ana[27] gpio_ana[28] gpio_ana[29] gpio_ana[30]
+ gpio_ana[31] gpio_ana[32] gpio_ana[33] gpio_ana[34] gpio_ana[35] gpio_ana[36] gpio_ana[37]
+ gpio_ana[38] gpio_ana[39] gpio_ana[40] gpio_ana[41] gpio_ana[42] gpio_ana[43] gpio_loopback_zero[0]
+ gpio_loopback_one[0] gpio_loopback_zero[1] gpio_loopback_one[1] gpio_loopback_zero[2]
+ gpio_loopback_one[2] gpio_loopback_one[3] gpio_loopback_zero[3] gpio_loopback_zero[4]
+ gpio_loopback_one[4] gpio_loopback_one[5] gpio_loopback_zero[5] gpio_loopback_zero[6]
+ gpio_loopback_one[6] gpio_loopback_one[7] gpio_loopback_zero[7] gpio_loopback_zero[8]
+ gpio_loopback_one[8] gpio_loopback_one[9] gpio_loopback_zero[9] gpio_loopback_zero[10]
+ gpio_loopback_one[10] gpio_loopback_one[11] gpio_loopback_zero[11] gpio_loopback_zero[12]
+ gpio_loopback_one[12] gpio_loopback_one[13] gpio_loopback_zero[14] gpio_loopback_one[14]
+ gpio_loopback_one[15] gpio_loopback_zero[15] gpio_loopback_zero[16] gpio_loopback_one[16]
+ gpio_loopback_one[17] gpio_loopback_zero[17] gpio_loopback_zero[18] gpio_loopback_one[18]
+ gpio_loopback_one[19] gpio_loopback_zero[19] gpio_loopback_zero[20] gpio_loopback_one[20]
+ gpio_loopback_one[21] gpio_loopback_zero[21] gpio_loopback_zero[22] gpio_loopback_one[22]
+ gpio_loopback_one[23] gpio_loopback_zero[23] gpio_loopback_zero[24] gpio_loopback_one[24]
+ gpio_loopback_one[25] gpio_loopback_zero[25] gpio_loopback_zero[26] gpio_loopback_one[26]
+ gpio_loopback_one[27] gpio_loopback_zero[27] gpio_loopback_zero[28] gpio_loopback_one[28]
+ gpio_loopback_one[29] gpio_loopback_zero[29] gpio_loopback_zero[30] gpio_loopback_one[30]
+ gpio_loopback_one[31] gpio_loopback_zero[31] gpio_loopback_zero[32] gpio_loopback_one[32]
+ gpio_loopback_one[33] gpio_loopback_zero[33] gpio_loopback_zero[34] gpio_loopback_one[34]
+ gpio_loopback_one[35] gpio_loopback_zero[35] gpio_loopback_zero[36] gpio_loopback_one[36]
+ gpio_loopback_one[37] gpio_loopback_zero[37] gpio_loopback_zero[38] gpio_loopback_one[38]
+ gpio_loopback_one[39] gpio_loopback_zero[39] gpio_loopback_zero[40] gpio_loopback_one[40]
+ gpio_loopback_one[41] gpio_loopback_zero[41] gpio_loopback_zero[42] gpio_loopback_one[42]
+ gpio_loopback_one[43] gpio_loopback_zero[43] resetb_pullup resetb_pulldown resetb_loopback_one
+ resetb_loopback_zero por_h porb_h porb_l mask_rev[0] mask_rev[1] mask_rev[2] mask_rev[3]
+ mask_rev[4] mask_rev[5] mask_rev[6] mask_rev[7] mask_rev[8] mask_rev[9] mask_rev[10]
+ mask_rev[11] mask_rev[12] mask_rev[13] mask_rev[14] mask_rev[15] mask_rev[16] mask_rev[17]
+ mask_rev[18] mask_rev[19] mask_rev[20] mask_rev[21] mask_rev[22] mask_rev[23] mask_rev[24]
+ mask_rev[25] mask_rev[26] mask_rev[27] mask_rev[28] mask_rev[29] mask_rev[30] mask_rev[31]
+ vssio vssd vddio vccd openframe_user_project_0/vert_connects_gpio_disabled_20/m2_32_13800#
+ openframe_user_project_0/vert_connects_gpio_disabled_18/m2_32_15194# openframe_user_project_0/vert_connects_gpio_disabled_18/m2_32_13800#
+ openframe_user_project_0/vert_connects_gpio_disabled_23/m2_32_13589# openframe_user_project_0/vert_connects_gpio_disabled_11/m2_32_2132#
+ openframe_user_project_0/vert_connects_gpio_disabled_8/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_13/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_13/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_16/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_12/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_9/m2_32_2132#
+ openframe_user_project_0/vert_connects_gpio_disabled_7/m2_32_14444# openframe_user_project_0/vert_connects_gpio_disabled_25/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_11/m2_32_13589# openframe_user_project_0/vert_connects_gpio_disabled_2/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_13/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_20/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_18/m2_32_14302# openframe_user_project_0/vert_connects_gpio_disabled_24/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_14/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_13/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_7/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_7/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_17/m2_32_14673# openframe_user_project_0/vert_connects_gpio_disabled_2/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_2/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_15/m2_32_2132#
+ openframe_user_project_0/vert_connects_gpio_disabled_12/m2_32_14673# openframe_user_project_0/vert_connects_gpio_disabled_5/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_16/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_0/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_24/m2_32_14444# openframe_user_project_0/vert_connects_gpio_disabled_7/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_17/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_17/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_2/m2_32_14302# openframe_user_project_0/vert_connects_gpio_disabled_6/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_18/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_12/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_1/m2_32_14673# openframe_user_project_0/vert_connects_gpio_disabled_24/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_24/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_19/m2_32_2132#
+ openframe_user_project_0/vert_connects_gpio_disabled_27/m2_32_13589# openframe_user_project_0/vert_connects_gpio_disabled_17/m2_32_13800#
+ openframe_user_project_0/vert_connects_gpio_disabled_17/m2_32_15194# openframe_user_project_0/vert_connects_gpio_disabled_22/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_12/m2_32_15194# openframe_user_project_0/vert_connects_gpio_disabled_12/m2_32_13800#
+ openframe_user_project_0/vert_connects_gpio_disabled_15/m2_32_13589# openframe_user_project_0/vert_connects_gpio_disabled_6/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_24/m2_32_14302# openframe_user_project_0/vert_connects_gpio_disabled_28/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_10/m2_32_13589# openframe_user_project_0/vert_connects_gpio_disabled_1/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_17/m2_32_14302# openframe_user_project_0/vert_connects_gpio_disabled_23/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_12/m2_32_14302# openframe_user_project_0/vert_connects_gpio_disabled_6/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_6/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_16/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_9/m2_32_13589# openframe_user_project_0/vert_connects_gpio_disabled_1/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_1/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_11/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_4/m2_32_13589# openframe_user_project_0/vert_connects_gpio_disabled_28/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_23/m2_32_14444# openframe_user_project_0/vert_connects_gpio_disabled_6/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_16/m2_32_14444# openframe_user_project_0/vert_connects_gpio_disabled_1/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_5/m2_32_14673# openframe_user_project_0/vert_connects_gpio_disabled_28/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_28/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_11/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_0/m2_32_14673# openframe_user_project_0/vert_connects_gpio_disabled_23/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_23/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_26/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_16/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_16/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_21/m2_32_13589# openframe_user_project_0/vert_connects_gpio_disabled_19/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_11/m2_32_15194# openframe_user_project_0/vert_connects_gpio_disabled_11/m2_32_13800#
+ gpio_drive1[19] openframe_user_project_0/vert_connects_gpio_disabled_28/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_14/m2_32_13589# openframe_user_project_0/vert_connects_gpio_disabled_5/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_23/m2_32_14302# openframe_user_project_0/vert_connects_gpio_disabled_27/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_0/m2_32_14444# openframe_user_project_0/vert_connects_gpio_disabled_16/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_22/m2_32_14673# openframe_user_project_0/vert_connects_gpio_disabled_11/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_5/m2_32_15194# openframe_user_project_0/vert_connects_gpio_disabled_15/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_5/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_8/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_0/m2_32_15194# openframe_user_project_0/vert_connects_gpio_disabled_0/m2_32_13800#
+ openframe_user_project_0/vert_connects_gpio_disabled_10/m2_32_14673# openframe_user_project_0/vert_connects_gpio_disabled_3/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_27/m2_32_14444# openframe_user_project_0/vert_connects_gpio_disabled_22/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_5/m2_32_14302# openframe_user_project_0/vert_connects_gpio_disabled_9/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_15/m2_32_14444# openframe_user_project_0/vert_connects_gpio_disabled_0/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_4/m2_32_14673# openframe_user_project_0/vert_connects_gpio_disabled_27/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_27/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_10/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_20/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_22/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_22/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_20/m2_32_1986#
+ openframe_user_project_0/vert_connects_gpio_disabled_25/m2_32_13589# openframe_user_project_0/vert_connects_gpio_disabled_15/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_21/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_15/m2_32_13800#
+ openframe_user_project_0/vert_connects_gpio_disabled_21/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_20/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_18/m2_32_13589# openframe_user_project_0/vert_connects_gpio_disabled_9/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_10/m2_32_15194# openframe_user_project_0/vert_connects_gpio_disabled_10/m2_32_13800#
+ openframe_user_project_0/vert_connects_gpio_disabled_27/m2_32_14302# openframe_user_project_0/vert_connects_gpio_disabled_22/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_0/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_22/m2_32_1986#
+ openframe_user_project_0/vert_connects_gpio_disabled_0/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_13/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_4/m2_32_14444# openframe_user_project_0/vert_connects_gpio_disabled_22/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_23/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_26/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_1/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_23/m2_32_1986#
+ openframe_user_project_0/vert_connects_gpio_disabled_1/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_15/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_21/m2_32_14673# openframe_user_project_0/vert_connects_gpio_disabled_9/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_19/m2_32_14673# openframe_user_project_0/vert_connects_gpio_disabled_9/m2_32_13800#
+ openframe_user_project_0/vert_connects_gpio_disabled_24/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_2/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_24/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_2/m2_32_1986#
+ openframe_user_project_0/vert_connects_gpio_disabled_10/m2_32_14302# openframe_user_project_0/vert_connects_gpio_disabled_4/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_4/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_14/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_25/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_7/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_3/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_25/m2_32_1986#
+ openframe_user_project_0/vert_connects_gpio_disabled_3/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_2/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_26/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_26/m2_32_1986#
+ openframe_user_project_0/vert_connects_gpio_disabled_4/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_4/m2_32_1986#
+ openframe_user_project_0/vert_connects_gpio_disabled_26/m2_32_14444# openframe_user_project_0/vert_connects_gpio_disabled_9/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_27/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_21/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_19/m2_32_14444# openframe_user_project_0/vert_connects_gpio_disabled_5/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_27/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_4/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_5/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_8/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_14/m2_32_14444# openframe_user_project_0/vert_connects_gpio_disabled_28/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_6/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_28/m2_32_1986#
+ openframe_user_project_0/vert_connects_gpio_disabled_3/m2_32_14673# openframe_user_project_0/vert_connects_gpio_disabled_6/m2_32_1986#
+ openframe_user_project_0/vert_connects_gpio_disabled_26/m2_32_15194# openframe_user_project_0/vert_connects_gpio_disabled_26/m2_32_13800#
+ openframe_user_project_0/vert_connects_gpio_disabled_20/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_10/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_21/m2_32_15194# openframe_user_project_0/vert_connects_gpio_disabled_7/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_21/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_10/m2_32_1986#
+ openframe_user_project_0/vert_connects_gpio_disabled_7/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_19/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_19/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_24/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_21/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_11/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_14/m2_32_15194# openframe_user_project_0/vert_connects_gpio_disabled_8/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_14/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_11/m2_32_1986#
+ openframe_user_project_0/vert_connects_gpio_disabled_8/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_17/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_22/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_8/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_0/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_9/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_26/m2_32_14302# openframe_user_project_0/vert_connects_gpio_disabled_12/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_12/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_9/m2_32_1986#
+ openframe_user_project_0/vert_connects_gpio_disabled_12/m2_32_13589# openframe_user_project_0/vert_connects_gpio_disabled_3/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_23/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_1/m2_32_2132#
+ openframe_user_project_0/vert_connects_gpio_disabled_21/m2_32_14302# openframe_user_project_0/vert_connects_gpio_disabled_19/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_13/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_25/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_13/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_24/m2_32_2132#
+ openframe_user_project_0/vert_connects_gpio_disabled_14/m2_32_14302# openframe_user_project_0/vert_connects_gpio_disabled_20/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_2/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_8/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_8/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_18/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_14/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_14/m2_32_1986#
+ openframe_user_project_0/vert_connects_gpio_disabled_3/m2_32_15194# openframe_user_project_0/vert_connects_gpio_disabled_25/m2_32_2132#
+ openframe_user_project_0/vert_connects_gpio_disabled_3/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_3/m2_32_2132#
+ gpio_loopback_zero[13] openframe_user_project_0/vert_connects_gpio_disabled_13/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_15/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_15/m2_32_1986#
+ openframe_user_project_0/vert_connects_gpio_disabled_6/m2_32_13589# openframe_user_project_0/vert_connects_gpio_disabled_26/m2_32_2132#
+ openframe_user_project_0/vert_connects_gpio_disabled_4/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_1/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_16/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_16/m2_32_1986#
+ openframe_user_project_0/vert_connects_gpio_disabled_25/m2_32_14444# openframe_user_project_0/vert_connects_gpio_disabled_8/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_27/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_5/m2_32_2132#
+ openframe_user_project_0/vert_connects_gpio_disabled_17/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_20/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_17/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_18/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_3/m2_32_14302# openframe_user_project_0/vert_connects_gpio_disabled_7/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_28/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_6/m2_32_2132#
+ openframe_user_project_0/vert_connects_gpio_disabled_13/m2_32_14444# openframe_user_project_0/vert_connects_gpio_disabled_18/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_18/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_2/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_25/m2_32_15194# openframe_user_project_0/vert_connects_gpio_disabled_25/m2_32_13800#
+ openframe_user_project_0/vert_connects_gpio_disabled_10/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_7/m2_32_2132#
+ openframe_user_project_0/vert_connects_gpio_disabled_28/m2_32_13589# openframe_user_project_0/vert_connects_gpio_disabled_19/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_20/m2_32_15194# openframe_user_project_0/vert_connects_gpio_disabled_19/m2_32_1986#
Xopenframe_user_project_0 gpio_in[38] gpio_in[40] gpio_oe[40] gpio_in[39] gpio_oe[39]
+ gpio_in[41] gpio_out[41] gpio_ie[41] gpio_oe[41] gpio_in[42] gpio_out[42] gpio_ie[42]
+ gpio_oe[42] gpio_drive0[38] gpio_drive1[38] gpio_in[43] gpio_ie[38] gpio_out[38]
+ gpio_oe[38] gpio_pulldown[38] gpio_pullup[38] gpio_schmitt[38] gpio_slew[38] gpio_schmitt[42]
+ gpio_pullup[42] gpio_drive0[42] gpio_drive1[42] gpio_pulldown[42] gpio_slew[42]
+ gpio_schmitt[41] gpio_pullup[41] gpio_drive0[41] gpio_drive1[41] gpio_pulldown[41]
+ gpio_slew[41] gpio_schmitt[40] gpio_pullup[40] gpio_drive0[40] gpio_drive1[40] gpio_pulldown[40]
+ gpio_ie[40] gpio_slew[40] gpio_out[40] gpio_schmitt[39] gpio_pullup[39] gpio_drive0[39]
+ gpio_drive1[39] gpio_pulldown[39] gpio_ie[39] gpio_slew[39] gpio_out[39] gpio_out[43]
+ gpio_slew[43] gpio_ie[43] gpio_pulldown[43] gpio_drive1[43] gpio_drive0[43] gpio_pullup[43]
+ gpio_schmitt[43] gpio_oe[43] gpio_drive0[30] gpio_drive0[0] gpio_drive0[5] gpio_drive1[5]
+ gpio_drive0[6] gpio_drive1[6] gpio_drive0[7] gpio_drive1[7] gpio_drive0[8] gpio_drive1[8]
+ gpio_drive0[9] gpio_drive1[9] gpio_drive1[0] gpio_drive0[10] gpio_drive1[10] gpio_drive0[11]
+ gpio_drive1[11] gpio_drive0[12] gpio_drive1[12] gpio_drive0[13] gpio_drive1[13]
+ gpio_drive0[14] gpio_drive1[14] gpio_drive0[1] gpio_drive0[15] gpio_drive0[16] gpio_drive1[16]
+ gpio_drive0[17] gpio_drive1[17] gpio_drive0[18] gpio_drive1[18] gpio_drive0[19]
+ gpio_drive1[19] gpio_drive1[1] gpio_drive0[20] gpio_drive1[20] gpio_drive0[21] gpio_drive1[21]
+ gpio_drive0[22] gpio_drive1[22] gpio_drive0[23] gpio_drive1[23] gpio_drive0[24]
+ gpio_drive1[24] gpio_drive0[2] gpio_drive1[25] gpio_drive0[25] gpio_drive0[26] gpio_drive1[26]
+ gpio_drive0[27] gpio_drive1[27] gpio_drive0[28] gpio_drive1[28] gpio_drive0[29]
+ gpio_drive1[29] gpio_drive1[2] gpio_drive1[30] gpio_drive0[31] gpio_drive1[31] gpio_drive0[32]
+ gpio_drive1[32] gpio_drive0[33] gpio_drive1[33] gpio_drive0[34] gpio_drive1[34]
+ gpio_drive0[3] gpio_drive0[35] gpio_drive1[35] gpio_drive0[36] gpio_drive1[36] gpio_drive0[37]
+ gpio_drive1[37] gpio_drive1[3] gpio_drive0[4] gpio_drive1[4] gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[34] gpio_in[35] gpio_in[36]
+ gpio_in[37] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_ie[0] gpio_ie[10] gpio_ie[11] gpio_ie[12] gpio_ie[13] gpio_ie[14] gpio_ie[15]
+ gpio_ie[16] gpio_ie[17] gpio_ie[18] gpio_ie[19] gpio_ie[1] gpio_ie[20] gpio_ie[21]
+ gpio_ie[22] gpio_ie[23] gpio_ie[24] gpio_ie[25] gpio_ie[26] gpio_ie[27] gpio_ie[28]
+ gpio_ie[29] gpio_ie[2] gpio_ie[30] gpio_ie[31] gpio_ie[32] gpio_ie[33] gpio_ie[34]
+ gpio_ie[35] gpio_ie[36] gpio_ie[37] gpio_ie[3] gpio_ie[4] gpio_ie[5] gpio_ie[6]
+ gpio_ie[7] gpio_ie[8] gpio_ie[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[34] gpio_out[35] gpio_out[36] gpio_out[37] gpio_out[3]
+ gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] gpio_oe[0]
+ gpio_oe[10] gpio_oe[11] gpio_oe[12] gpio_oe[13] gpio_oe[14] gpio_oe[15] gpio_oe[16]
+ gpio_oe[17] gpio_oe[18] gpio_oe[19] gpio_oe[1] gpio_oe[20] gpio_oe[21] gpio_oe[22]
+ gpio_oe[23] gpio_oe[24] gpio_oe[25] gpio_oe[26] gpio_oe[27] gpio_oe[28] gpio_oe[29]
+ gpio_oe[2] gpio_oe[30] gpio_oe[31] gpio_oe[32] gpio_oe[33] gpio_oe[34] gpio_oe[35]
+ gpio_oe[36] gpio_oe[37] gpio_oe[3] gpio_oe[4] gpio_oe[5] gpio_oe[6] gpio_oe[7] gpio_oe[8]
+ gpio_oe[9] gpio_pulldown[0] gpio_pulldown[10] gpio_pulldown[11] gpio_pulldown[12]
+ gpio_pulldown[13] gpio_pulldown[14] gpio_pulldown[15] gpio_pulldown[16] gpio_pulldown[17]
+ gpio_pulldown[18] gpio_pulldown[19] gpio_pulldown[1] gpio_pulldown[20] gpio_pulldown[21]
+ gpio_pulldown[22] gpio_pulldown[23] gpio_pulldown[24] gpio_pulldown[25] gpio_pulldown[26]
+ gpio_pulldown[27] gpio_pulldown[28] gpio_pulldown[29] gpio_pulldown[2] gpio_pulldown[30]
+ gpio_pulldown[31] gpio_pulldown[32] gpio_pulldown[33] gpio_pulldown[34] gpio_pulldown[35]
+ gpio_pulldown[36] gpio_pulldown[37] gpio_pulldown[3] gpio_pulldown[4] gpio_pulldown[5]
+ gpio_pulldown[6] gpio_pulldown[7] gpio_pulldown[8] gpio_pulldown[9] gpio_pullup[0]
+ gpio_pullup[10] gpio_pullup[11] gpio_pullup[12] gpio_pullup[13] gpio_pullup[14]
+ gpio_pullup[15] gpio_pullup[16] gpio_pullup[17] gpio_pullup[18] gpio_pullup[19]
+ gpio_pullup[1] gpio_pullup[20] gpio_pullup[21] gpio_pullup[22] gpio_pullup[23] gpio_pullup[24]
+ gpio_pullup[25] gpio_pullup[26] gpio_pullup[27] gpio_pullup[28] gpio_pullup[29]
+ gpio_pullup[2] gpio_pullup[30] gpio_pullup[31] gpio_pullup[32] gpio_pullup[33] gpio_pullup[34]
+ gpio_pullup[35] gpio_pullup[36] gpio_pullup[37] gpio_pullup[3] gpio_pullup[4] gpio_pullup[5]
+ gpio_pullup[6] gpio_pullup[7] gpio_pullup[8] gpio_pullup[9] gpio_schmitt[0] gpio_schmitt[10]
+ gpio_schmitt[11] gpio_schmitt[12] gpio_schmitt[13] gpio_schmitt[14] gpio_schmitt[15]
+ gpio_schmitt[16] gpio_schmitt[17] gpio_schmitt[18] gpio_schmitt[19] gpio_schmitt[1]
+ gpio_schmitt[20] gpio_schmitt[21] gpio_schmitt[22] gpio_schmitt[23] gpio_schmitt[24]
+ gpio_schmitt[25] gpio_schmitt[26] gpio_schmitt[27] gpio_schmitt[28] gpio_schmitt[29]
+ gpio_schmitt[2] gpio_schmitt[30] gpio_schmitt[31] gpio_schmitt[32] gpio_schmitt[33]
+ gpio_schmitt[34] gpio_schmitt[35] gpio_schmitt[36] gpio_schmitt[37] gpio_schmitt[3]
+ gpio_schmitt[4] gpio_schmitt[5] gpio_schmitt[6] gpio_schmitt[7] gpio_schmitt[8]
+ gpio_schmitt[9] gpio_slew[0] gpio_slew[10] gpio_slew[11] gpio_slew[12] gpio_slew[13]
+ gpio_slew[14] gpio_slew[15] gpio_slew[16] gpio_slew[17] gpio_slew[18] gpio_slew[19]
+ gpio_slew[1] gpio_slew[20] gpio_slew[21] gpio_slew[22] gpio_slew[23] gpio_slew[24]
+ gpio_slew[25] gpio_slew[26] gpio_slew[27] gpio_slew[28] gpio_slew[29] gpio_slew[2]
+ gpio_slew[30] gpio_slew[31] gpio_slew[32] gpio_slew[33] gpio_slew[34] gpio_slew[35]
+ gpio_slew[36] gpio_slew[37] gpio_slew[3] gpio_slew[4] gpio_slew[5] gpio_slew[6]
+ gpio_slew[7] gpio_slew[8] gpio_slew[9] resetb_core gpio_ana[0] gpio_ana[1] gpio_ana[2]
+ gpio_ana[3] gpio_ana[4] gpio_ana[5] gpio_ana[6] gpio_ana[7] gpio_ana[8] gpio_ana[9]
+ gpio_ana[10] gpio_ana[11] gpio_ana[12] gpio_ana[13] gpio_ana[14] gpio_ana[15] gpio_ana[16]
+ gpio_ana[17] gpio_ana[18] gpio_ana[19] gpio_ana[20] gpio_ana[21] gpio_ana[22] gpio_ana[23]
+ gpio_ana[24] gpio_ana[25] gpio_ana[26] gpio_ana[27] gpio_ana[28] gpio_ana[29] gpio_ana[30]
+ gpio_ana[31] gpio_ana[32] gpio_ana[33] gpio_ana[34] gpio_ana[35] gpio_ana[36] gpio_ana[37]
+ gpio_ana[38] gpio_ana[39] gpio_ana[40] gpio_ana[41] gpio_ana[42] gpio_ana[43] gpio_loopback_zero[0]
+ gpio_loopback_one[0] gpio_loopback_zero[1] gpio_loopback_one[1] gpio_loopback_zero[2]
+ gpio_loopback_one[2] gpio_loopback_one[3] gpio_loopback_zero[3] gpio_loopback_zero[4]
+ gpio_loopback_one[4] gpio_loopback_one[5] gpio_loopback_zero[5] gpio_loopback_zero[6]
+ gpio_loopback_one[6] gpio_loopback_one[7] gpio_loopback_zero[7] gpio_loopback_zero[8]
+ gpio_loopback_one[8] gpio_loopback_one[9] gpio_loopback_zero[9] gpio_loopback_zero[10]
+ gpio_loopback_one[10] gpio_loopback_one[11] gpio_loopback_zero[11] gpio_loopback_zero[12]
+ gpio_loopback_one[12] gpio_loopback_one[13] gpio_loopback_zero[13] gpio_loopback_zero[14]
+ gpio_loopback_one[14] gpio_loopback_one[15] gpio_loopback_zero[15] gpio_loopback_zero[16]
+ gpio_loopback_one[16] gpio_loopback_one[17] gpio_loopback_zero[17] gpio_loopback_zero[18]
+ gpio_loopback_one[18] gpio_loopback_one[19] gpio_loopback_zero[19] gpio_loopback_zero[20]
+ gpio_loopback_one[20] gpio_loopback_one[21] gpio_loopback_zero[21] gpio_loopback_zero[22]
+ gpio_loopback_one[22] gpio_loopback_one[23] gpio_loopback_zero[23] gpio_loopback_zero[24]
+ gpio_loopback_one[24] gpio_loopback_one[25] gpio_loopback_zero[25] gpio_loopback_zero[26]
+ gpio_loopback_one[26] gpio_loopback_one[27] gpio_loopback_zero[27] gpio_loopback_zero[28]
+ gpio_loopback_one[28] gpio_loopback_one[29] gpio_loopback_zero[29] gpio_loopback_zero[30]
+ gpio_loopback_one[30] gpio_loopback_one[31] gpio_loopback_zero[31] gpio_loopback_zero[32]
+ gpio_loopback_one[32] gpio_loopback_one[33] gpio_loopback_zero[33] gpio_loopback_zero[34]
+ gpio_loopback_one[34] gpio_loopback_one[35] gpio_loopback_zero[35] gpio_loopback_zero[36]
+ gpio_loopback_one[36] gpio_loopback_one[37] gpio_loopback_zero[37] gpio_loopback_zero[38]
+ gpio_loopback_one[38] gpio_loopback_one[39] gpio_loopback_zero[39] gpio_loopback_zero[40]
+ gpio_loopback_one[40] gpio_loopback_one[41] gpio_loopback_zero[41] gpio_loopback_zero[42]
+ gpio_loopback_one[42] gpio_loopback_one[43] gpio_loopback_zero[43] resetb_pullup
+ resetb_pulldown resetb_loopback_one resetb_loopback_zero por_h porb_h porb_l mask_rev[0]
+ mask_rev[1] mask_rev[2] mask_rev[3] mask_rev[4] mask_rev[5] mask_rev[6] mask_rev[7]
+ mask_rev[8] mask_rev[9] mask_rev[10] mask_rev[11] mask_rev[12] mask_rev[13] mask_rev[14]
+ mask_rev[15] mask_rev[16] mask_rev[17] mask_rev[18] mask_rev[19] mask_rev[20] mask_rev[21]
+ mask_rev[22] mask_rev[23] mask_rev[24] mask_rev[25] mask_rev[26] mask_rev[27] mask_rev[28]
+ mask_rev[29] mask_rev[30] mask_rev[31] vssio vssd vddio vccd openframe_user_project_0/vert_connects_gpio_disabled_15/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_27/m2_32_15194# openframe_user_project_0/vert_connects_gpio_disabled_27/m2_32_13800#
+ openframe_user_project_0/vert_connects_gpio_disabled_10/m2_32_14444# openframe_user_project_0/vert_connects_gpio_disabled_22/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_22/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_25/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_15/m2_32_15194# openframe_user_project_0/vert_connects_gpio_disabled_5/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_15/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_20/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_18/m2_32_13589# openframe_user_project_0/vert_connects_gpio_disabled_10/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_0/m2_32_14444# openframe_user_project_0/vert_connects_gpio_disabled_10/m2_32_13800#
+ openframe_user_project_0/vert_connects_gpio_disabled_27/m2_32_14302# openframe_user_project_0/vert_connects_gpio_disabled_13/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_22/m2_32_14302# openframe_user_project_0/vert_connects_gpio_disabled_26/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_5/m2_32_15194# openframe_user_project_0/vert_connects_gpio_disabled_5/m2_32_13800#
+ openframe_user_project_0/vert_connects_gpio_disabled_8/m2_32_13589# openframe_user_project_0/vert_connects_gpio_disabled_15/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_21/m2_32_14673# openframe_user_project_0/vert_connects_gpio_disabled_0/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_0/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_19/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_3/m2_32_13589# openframe_user_project_0/vert_connects_gpio_disabled_10/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_14/m2_32_14673# openframe_user_project_0/vert_connects_gpio_disabled_5/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_9/m2_32_14673# openframe_user_project_0/vert_connects_gpio_disabled_26/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_0/m2_32_14302# openframe_user_project_0/vert_connects_gpio_disabled_4/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_21/m2_32_14444# openframe_user_project_0/vert_connects_gpio_disabled_19/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_20/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_20/m2_32_1986#
+ openframe_user_project_0/vert_connects_gpio_disabled_14/m2_32_14444# openframe_user_project_0/vert_connects_gpio_disabled_26/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_26/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_21/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_21/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_21/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_21/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_19/m2_32_13800#
+ openframe_user_project_0/vert_connects_gpio_disabled_9/m2_32_14444# openframe_user_project_0/vert_connects_gpio_disabled_19/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_22/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_24/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_22/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_14/m2_32_13800#
+ openframe_user_project_0/vert_connects_gpio_disabled_14/m2_32_15194# openframe_user_project_0/vert_connects_gpio_disabled_4/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_23/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_17/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_23/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_26/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_12/m2_32_13589# openframe_user_project_0/vert_connects_gpio_disabled_9/m2_32_13800#
+ openframe_user_project_0/vert_connects_gpio_disabled_9/m2_32_15194# openframe_user_project_0/vert_connects_gpio_disabled_24/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_24/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_21/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_19/m2_32_14302# openframe_user_project_0/vert_connects_gpio_disabled_25/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_4/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_4/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_25/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_7/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_25/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_14/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_20/m2_32_14673# openframe_user_project_0/vert_connects_gpio_disabled_18/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_2/m2_32_13589# openframe_user_project_0/vert_connects_gpio_disabled_26/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_13/m2_32_14673# openframe_user_project_0/vert_connects_gpio_disabled_26/m2_32_1986#
+ openframe_user_project_0/vert_connects_gpio_disabled_9/m2_32_14302# openframe_user_project_0/vert_connects_gpio_disabled_0/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_0/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_27/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_27/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_4/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_8/m2_32_14673# openframe_user_project_0/vert_connects_gpio_disabled_25/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_1/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_28/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_1/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_28/m2_32_1986#
+ openframe_user_project_0/vert_connects_gpio_disabled_3/m2_32_14673# openframe_user_project_0/vert_connects_gpio_disabled_20/m2_32_14444#
+ gpio_drive1[15] openframe_user_project_0/vert_connects_gpio_disabled_20/m2_32_2132#
+ openframe_user_project_0/vert_connects_gpio_disabled_18/m2_32_14444# openframe_user_project_0/vert_connects_gpio_disabled_2/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_10/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_2/m2_32_1986#
+ openframe_user_project_0/vert_connects_gpio_disabled_10/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_13/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_21/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_25/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_3/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_25/m2_32_13800#
+ openframe_user_project_0/vert_connects_gpio_disabled_3/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_11/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_11/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_28/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_22/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_20/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_20/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_8/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_18/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_18/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_4/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_12/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_4/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_23/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_12/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_13/m2_32_13800#
+ openframe_user_project_0/vert_connects_gpio_disabled_13/m2_32_15194# openframe_user_project_0/vert_connects_gpio_disabled_3/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_23/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_5/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_5/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_13/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_16/m2_32_13589# openframe_user_project_0/vert_connects_gpio_disabled_13/m2_32_1986#
+ openframe_user_project_0/vert_connects_gpio_disabled_25/m2_32_14302# openframe_user_project_0/vert_connects_gpio_disabled_24/m2_32_2132#
+ openframe_user_project_0/vert_connects_gpio_disabled_8/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_6/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_8/m2_32_15194# openframe_user_project_0/vert_connects_gpio_disabled_11/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_14/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_6/m2_32_1986#
+ openframe_user_project_0/vert_connects_gpio_disabled_14/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_20/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_18/m2_32_14302# openframe_user_project_0/vert_connects_gpio_disabled_24/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_3/m2_32_15194# openframe_user_project_0/vert_connects_gpio_disabled_25/m2_32_2132#
+ openframe_user_project_0/vert_connects_gpio_disabled_3/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_7/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_7/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_15/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_15/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_6/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_13/m2_32_14302# openframe_user_project_0/vert_connects_gpio_disabled_17/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_26/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_8/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_1/m2_32_13589# openframe_user_project_0/vert_connects_gpio_disabled_8/m2_32_1986#
+ openframe_user_project_0/vert_connects_gpio_disabled_16/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_12/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_16/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_8/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_0/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_27/m2_32_2132#
+ openframe_user_project_0/vert_connects_gpio_disabled_9/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_9/m2_32_1986#
+ openframe_user_project_0/vert_connects_gpio_disabled_17/m2_32_1840# openframe_user_project_0/vert_connects_gpio_disabled_17/m2_32_1986#
+ openframe_user_project_0/vert_connects_gpio_disabled_3/m2_32_14302# openframe_user_project_0/vert_connects_gpio_disabled_7/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_1/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_28/m2_32_2132#
+ openframe_user_project_0/vert_connects_gpio_disabled_24/m2_32_14444# openframe_user_project_0/vert_connects_gpio_disabled_18/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_18/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_2/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_2/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_10/m2_32_2132#
+ openframe_user_project_0/vert_connects_gpio_disabled_17/m2_32_14444# openframe_user_project_0/vert_connects_gpio_disabled_19/m2_32_1840#
+ openframe_user_project_0/vert_connects_gpio_disabled_19/m2_32_1986# openframe_user_project_0/vert_connects_gpio_disabled_12/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_3/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_11/m2_32_2132#
+ openframe_user_project_0/vert_connects_gpio_disabled_24/m2_32_15194# openframe_user_project_0/vert_connects_gpio_disabled_24/m2_32_13800#
+ openframe_user_project_0/vert_connects_gpio_disabled_27/m2_32_13589# openframe_user_project_0/vert_connects_gpio_disabled_4/m2_32_2132#
+ openframe_user_project_0/vert_connects_gpio_disabled_12/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_7/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_17/m2_32_15194# openframe_user_project_0/vert_connects_gpio_disabled_17/m2_32_13800#
+ openframe_user_project_0/vert_connects_gpio_disabled_22/m2_32_13589# openframe_user_project_0/vert_connects_gpio_disabled_5/m2_32_2132#
+ openframe_user_project_0/vert_connects_gpio_disabled_2/m2_32_14444# openframe_user_project_0/vert_connects_gpio_disabled_12/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_12/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_13/m2_32_2132#
+ openframe_user_project_0/vert_connects_gpio_disabled_15/m2_32_13589# openframe_user_project_0/vert_connects_gpio_disabled_6/m2_32_2132#
+ openframe_user_project_0/vert_connects_gpio_disabled_24/m2_32_14302# openframe_user_project_0/vert_connects_gpio_disabled_14/m2_32_2132#
+ openframe_user_project_0/vert_connects_gpio_disabled_28/m2_32_14673# openframe_user_project_0/vert_connects_gpio_disabled_10/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_7/m2_32_15194# openframe_user_project_0/vert_connects_gpio_disabled_7/m2_32_13800#
+ openframe_user_project_0/vert_connects_gpio_disabled_7/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_17/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_23/m2_32_14673# openframe_user_project_0/vert_connects_gpio_disabled_2/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_15/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_2/m2_32_13800#
+ openframe_user_project_0/vert_connects_gpio_disabled_5/m2_32_13589# openframe_user_project_0/vert_connects_gpio_disabled_12/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_16/m2_32_14673# openframe_user_project_0/vert_connects_gpio_disabled_8/m2_32_2132#
+ openframe_user_project_0/vert_connects_gpio_disabled_16/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_0/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_11/m2_32_14673# openframe_user_project_0/vert_connects_gpio_disabled_9/m2_32_2132#
+ openframe_user_project_0/vert_connects_gpio_disabled_7/m2_32_14302# openframe_user_project_0/vert_connects_gpio_disabled_17/m2_32_2132#
+ openframe_user_project_0/vert_connects_gpio_disabled_28/m2_32_14444# openframe_user_project_0/vert_connects_gpio_disabled_2/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_6/m2_32_14673# openframe_user_project_0/vert_connects_gpio_disabled_18/m2_32_2132#
+ openframe_user_project_0/vert_connects_gpio_disabled_23/m2_32_14444# openframe_user_project_0/vert_connects_gpio_disabled_1/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_19/m2_32_2132# openframe_user_project_0/vert_connects_gpio_disabled_16/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_28/m2_32_15194# openframe_user_project_0/vert_connects_gpio_disabled_28/m2_32_13800#
+ openframe_user_project_0/vert_connects_gpio_disabled_11/m2_32_14444# openframe_user_project_0/vert_connects_gpio_disabled_23/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_23/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_26/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_16/m2_32_15194# openframe_user_project_0/vert_connects_gpio_disabled_16/m2_32_13800#
+ openframe_user_project_0/vert_connects_gpio_disabled_6/m2_32_14444# openframe_user_project_0/vert_connects_gpio_disabled_21/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_19/m2_32_13589# openframe_user_project_0/vert_connects_gpio_disabled_11/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_11/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_1/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_28/m2_32_14302# openframe_user_project_0/vert_connects_gpio_disabled_14/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_23/m2_32_14302# openframe_user_project_0/vert_connects_gpio_disabled_27/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_6/m2_32_15194# openframe_user_project_0/vert_connects_gpio_disabled_6/m2_32_13800#
+ openframe_user_project_0/vert_connects_gpio_disabled_9/m2_32_13589# openframe_user_project_0/vert_connects_gpio_disabled_16/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_22/m2_32_14673# openframe_user_project_0/vert_connects_gpio_disabled_1/m2_32_15194#
+ openframe_user_project_0/vert_connects_gpio_disabled_1/m2_32_13800# openframe_user_project_0/vert_connects_gpio_disabled_4/m2_32_13589#
+ openframe_user_project_0/vert_connects_gpio_disabled_11/m2_32_14302# openframe_user_project_0/vert_connects_gpio_disabled_15/m2_32_14673#
+ openframe_user_project_0/vert_connects_gpio_disabled_10/m2_32_14673# openframe_user_project_0/vert_connects_gpio_disabled_6/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_27/m2_32_14444# openframe_user_project_0/vert_connects_gpio_disabled_1/m2_32_14302#
+ openframe_user_project_0/vert_connects_gpio_disabled_5/m2_32_14673# openframe_user_project_0/vert_connects_gpio_disabled_22/m2_32_14444#
+ openframe_user_project_0/vert_connects_gpio_disabled_0/m2_32_14673# openframe_user_project
.ends

.subckt caravel_openframe vddio gpio[38] gpio[39] gpio[40] gpio[41] gpio[42] gpio[43]
+ gpio[0] gpio[10] gpio[11] gpio[12] gpio[13] gpio[14] gpio[15] gpio[16] gpio[17]
+ gpio[18] gpio[19] gpio[1] gpio[20] gpio[21] gpio[22] gpio[23] gpio[24] gpio[25]
+ gpio[26] gpio[27] gpio[28] gpio[29] gpio[2] gpio[30] gpio[31] gpio[32] gpio[33]
+ gpio[34] gpio[35] gpio[36] gpio[37] gpio[3] gpio[4] gpio[5] gpio[6] gpio[7] gpio[8]
+ gpio[9] resetb vssd vccd
Xpadframe padframe/gpio_in[38] gpio[39] padframe/gpio_in[39] padframe/gpio_drive2[38]
+ padframe/gpio_in[43] gpio[10] gpio[13] gpio[16] gpio[19] gpio[22] gpio[25] gpio[2]
+ gpio[30] gpio[32] gpio[33] gpio[35] gpio[36] padframe/gpio_drive0[0] padframe/gpio_drive0[5]
+ padframe/gpio_drive1[6] padframe/gpio_drive1[7] padframe/gpio_drive1[8] padframe/gpio_drive0[9]
+ padframe/gpio_drive1[9] padframe/gpio_drive0[10] padframe/gpio_drive0[11] padframe/gpio_drive0[12]
+ padframe/gpio_drive0[13] padframe/gpio_drive1[13] padframe/gpio_drive0[14] padframe/gpio_drive0[1]
+ padframe/gpio_drive0[15] padframe/gpio_drive0[16] padframe/gpio_drive0[17] padframe/gpio_drive0[18]
+ padframe/gpio_drive1[18] padframe/gpio_drive1[1] padframe/gpio_drive1[21] padframe/gpio_drive1[22]
+ padframe/gpio_drive0[23] padframe/gpio_drive1[23] padframe/gpio_drive0[24] padframe/gpio_drive1[24]
+ padframe/gpio_drive0[2] padframe/gpio_drive1[26] padframe/gpio_drive1[27] padframe/gpio_drive0[28]
+ padframe/gpio_drive1[28] padframe/gpio_drive0[29] padframe/gpio_drive1[29] padframe/gpio_drive1[2]
+ padframe/gpio_drive1[30] padframe/gpio_drive0[32] padframe/gpio_drive0[33] padframe/gpio_drive0[34]
+ padframe/gpio_drive0[3] padframe/gpio_drive0[35] padframe/gpio_drive1[35] padframe/gpio_drive0[36]
+ padframe/gpio_drive1[3] padframe/gpio_in[0] padframe/gpio_in[10] padframe/gpio_in[11]
+ padframe/gpio_in[12] padframe/gpio_in[13] padframe/gpio_in[14] padframe/gpio_in[15]
+ padframe/gpio_in[16] padframe/gpio_in[17] padframe/gpio_in[18] padframe/gpio_in[19]
+ padframe/gpio_in[1] padframe/gpio_in[25] padframe/gpio_in[26] padframe/gpio_in[27]
+ padframe/gpio_in[29] padframe/gpio_in[2] padframe/gpio_in[30] padframe/gpio_in[31]
+ padframe/gpio_in[32] padframe/gpio_in[33] padframe/gpio_in[34] padframe/gpio_in[35]
+ padframe/gpio_in[36] padframe/gpio_in[37] padframe/gpio_in[3] padframe/gpio_in[4]
+ padframe/gpio_in[5] padframe/gpio_in[7] padframe/gpio_in[8] padframe/gpio_in[9]
+ padframe/gpio_ie[10] padframe/gpio_ie[11] padframe/gpio_ie[12] padframe/gpio_ie[13]
+ padframe/gpio_ie[14] padframe/gpio_ie[24] padframe/gpio_ie[25] padframe/gpio_ie[28]
+ padframe/gpio_ie[29] padframe/gpio_ie[2] padframe/gpio_ie[30] padframe/gpio_ie[33]
+ padframe/gpio_ie[5] padframe/gpio_ie[6] padframe/gpio_ie[9] padframe/gpio_out[10]
+ padframe/gpio_out[11] padframe/gpio_out[13] padframe/gpio_out[14] padframe/gpio_out[17]
+ padframe/gpio_out[19] padframe/gpio_out[22] padframe/gpio_out[25] padframe/gpio_out[28]
+ padframe/gpio_out[30] padframe/gpio_out[32] padframe/gpio_out[33] padframe/gpio_out[34]
+ padframe/gpio_out[35] padframe/gpio_out[36] padframe/gpio_out[37] padframe/gpio_out[6]
+ padframe/gpio_out[9] padframe/gpio_oe[10] padframe/gpio_oe[12] padframe/gpio_oe[13]
+ padframe/gpio_oe[15] padframe/gpio_oe[16] padframe/gpio_oe[17] padframe/gpio_oe[18]
+ padframe/gpio_oe[19] padframe/gpio_oe[24] padframe/gpio_oe[27] padframe/gpio_oe[28]
+ padframe/gpio_oe[30] padframe/gpio_oe[31] padframe/gpio_oe[33] padframe/gpio_oe[34]
+ padframe/gpio_oe[35] padframe/gpio_oe[36] padframe/gpio_oe[8] padframe/gpio_pulldown[11]
+ padframe/gpio_pulldown[15] padframe/gpio_pulldown[1] padframe/gpio_pulldown[21]
+ padframe/gpio_pulldown[22] padframe/gpio_pulldown[24] padframe/gpio_pulldown[25]
+ padframe/gpio_pulldown[27] padframe/gpio_pulldown[28] padframe/gpio_pulldown[29]
+ padframe/gpio_pulldown[2] padframe/gpio_pulldown[33] padframe/gpio_pulldown[36]
+ padframe/gpio_pulldown[5] padframe/gpio_pulldown[8] padframe/gpio_pulldown[9] padframe/gpio_pullup[0]
+ padframe/gpio_pullup[10] padframe/gpio_pullup[11] padframe/gpio_pullup[12] padframe/gpio_pullup[13]
+ padframe/gpio_pullup[14] padframe/gpio_pullup[15] padframe/gpio_pullup[1] padframe/gpio_pullup[25]
+ padframe/gpio_pullup[26] padframe/gpio_pullup[28] padframe/gpio_pullup[29] padframe/gpio_pullup[30]
+ padframe/gpio_pullup[31] padframe/gpio_pullup[32] padframe/gpio_pullup[33] padframe/gpio_pullup[37]
+ padframe/gpio_pullup[3] padframe/gpio_pullup[4] padframe/gpio_pullup[6] padframe/gpio_pullup[7]
+ padframe/gpio_pullup[8] padframe/gpio_pullup[9] padframe/gpio_schmitt[11] padframe/gpio_schmitt[12]
+ padframe/gpio_schmitt[13] padframe/gpio_schmitt[14] padframe/gpio_schmitt[15] padframe/gpio_schmitt[1]
+ padframe/gpio_schmitt[20] padframe/gpio_schmitt[24] padframe/gpio_schmitt[26] padframe/gpio_schmitt[27]
+ padframe/gpio_schmitt[29] padframe/gpio_schmitt[2] padframe/gpio_schmitt[30] padframe/gpio_schmitt[31]
+ padframe/gpio_schmitt[32] padframe/gpio_schmitt[4] padframe/gpio_schmitt[5] padframe/gpio_schmitt[6]
+ padframe/gpio_schmitt[7] padframe/gpio_schmitt[8] padframe/gpio_schmitt[9] padframe/gpio_slew[0]
+ padframe/gpio_slew[15] padframe/gpio_slew[22] padframe/gpio_slew[24] padframe/gpio_slew[25]
+ padframe/gpio_slew[26] padframe/gpio_slew[27] padframe/gpio_slew[28] padframe/gpio_slew[29]
+ padframe/gpio_slew[2] padframe/gpio_slew[33] padframe/gpio_slew[36] padframe/gpio_slew[3]
+ padframe/gpio_slew[4] padframe/gpio_slew[5] padframe/gpio_slew[6] padframe/gpio_slew[7]
+ padframe/gpio_slew[8] padframe/gpio_slew[9] padframe/resetb_core padframe/gpio_ana[0]
+ padframe/gpio_ana[1] padframe/gpio_ana[2] padframe/gpio_ana[3] padframe/gpio_ana[4]
+ padframe/gpio_ana[5] padframe/gpio_ana[6] padframe/gpio_ana[7] padframe/gpio_ana[8]
+ padframe/gpio_ana[9] padframe/gpio_ana[10] padframe/gpio_ana[11] padframe/gpio_ana[12]
+ padframe/gpio_ana[13] padframe/gpio_ana[14] padframe/gpio_ana[18] padframe/gpio_ana[21]
+ padframe/gpio_ana[22] padframe/gpio_ana[23] padframe/gpio_ana[24] padframe/gpio_ana[25]
+ padframe/gpio_ana[26] padframe/gpio_ana[27] padframe/gpio_ana[28] padframe/gpio_ana[29]
+ padframe/gpio_ana[30] padframe/gpio_ana[31] padframe/gpio_ana[32] padframe/gpio_ana[33]
+ padframe/gpio_ana[34] padframe/gpio_ana[35] padframe/gpio_ana[36] padframe/gpio_ana[37]
+ padframe/gpio_ana[40] padframe/gpio_ana[41] padframe/gpio_ana[42] padframe/gpio_ana[43]
+ padframe/gpio_loopback_zero[0] padframe/gpio_loopback_one[0] padframe/gpio_loopback_zero[1]
+ padframe/gpio_loopback_one[1] padframe/gpio_loopback_zero[2] padframe/gpio_loopback_one[2]
+ padframe/gpio_loopback_one[3] padframe/gpio_loopback_zero[3] padframe/gpio_loopback_zero[4]
+ padframe/gpio_loopback_one[4] padframe/gpio_loopback_one[5] padframe/gpio_loopback_zero[5]
+ padframe/gpio_loopback_zero[6] padframe/gpio_loopback_one[6] padframe/gpio_loopback_one[7]
+ padframe/gpio_loopback_zero[7] padframe/gpio_loopback_zero[8] padframe/gpio_loopback_one[8]
+ padframe/gpio_loopback_one[9] padframe/gpio_loopback_zero[9] padframe/gpio_loopback_zero[10]
+ padframe/gpio_loopback_one[11] padframe/gpio_loopback_zero[11] padframe/gpio_loopback_zero[12]
+ padframe/gpio_loopback_one[12] padframe/gpio_loopback_one[13] padframe/gpio_loopback_zero[14]
+ padframe/gpio_loopback_one[14] padframe/gpio_loopback_one[15] padframe/gpio_loopback_zero[15]
+ padframe/gpio_loopback_zero[16] padframe/gpio_loopback_one[16] padframe/gpio_loopback_one[17]
+ padframe/gpio_loopback_zero[17] padframe/gpio_loopback_zero[18] padframe/gpio_loopback_one[18]
+ padframe/gpio_loopback_one[19] padframe/gpio_loopback_zero[19] padframe/gpio_loopback_zero[20]
+ padframe/gpio_loopback_one[20] padframe/gpio_loopback_one[21] padframe/gpio_loopback_zero[21]
+ padframe/gpio_loopback_one[22] padframe/gpio_loopback_one[23] padframe/gpio_loopback_zero[23]
+ padframe/gpio_loopback_zero[24] padframe/gpio_loopback_one[25] padframe/gpio_loopback_zero[25]
+ padframe/gpio_loopback_zero[26] padframe/gpio_loopback_one[26] padframe/gpio_loopback_one[27]
+ padframe/gpio_loopback_zero[27] padframe/gpio_loopback_zero[28] padframe/gpio_loopback_one[28]
+ padframe/gpio_loopback_one[29] padframe/gpio_loopback_zero[29] padframe/gpio_loopback_zero[30]
+ padframe/gpio_loopback_one[30] padframe/gpio_loopback_one[31] padframe/gpio_loopback_zero[31]
+ padframe/gpio_loopback_zero[32] padframe/gpio_loopback_one[32] padframe/gpio_loopback_zero[33]
+ padframe/gpio_loopback_zero[34] padframe/gpio_loopback_one[34] padframe/gpio_loopback_one[35]
+ padframe/gpio_loopback_zero[35] padframe/gpio_loopback_zero[36] padframe/gpio_loopback_one[36]
+ padframe/gpio_loopback_one[37] padframe/gpio_loopback_zero[37] padframe/gpio_loopback_zero[38]
+ padframe/gpio_loopback_zero[39] padframe/gpio_loopback_zero[40] padframe/gpio_loopback_one[40]
+ padframe/gpio_loopback_one[41] padframe/gpio_loopback_one[43] padframe/gpio_loopback_zero[43]
+ padframe/resetb_loopback_zero padframe/porb_h padframe/porb_l padframe/mask_rev[0]
+ padframe/mask_rev[1] padframe/mask_rev[2] padframe/mask_rev[3] padframe/mask_rev[4]
+ padframe/mask_rev[5] padframe/mask_rev[6] padframe/mask_rev[7] padframe/mask_rev[8]
+ padframe/mask_rev[9] padframe/mask_rev[20] padframe/mask_rev[21] padframe/mask_rev[22]
+ padframe/mask_rev[23] padframe/mask_rev[24] padframe/mask_rev[25] padframe/mask_rev[26]
+ padframe/gpio_drive0[30] padframe/gpio_drive0[42] padframe/gpio_drive1[42] padframe/gpio_pulldown[42]
+ padframe/gpio_pullup[41] padframe/gpio_drive0[41] padframe/gpio_drive1[41] padframe/gpio_slew[41]
+ padframe/gpio_schmitt[40] padframe/gpio_out[39] padframe/gpio_oe[43] padframe/gpio_slew[43]
+ padframe/gpio_ie[43] padframe/gpio_pulldown[43] padframe/gpio_drive1[43] padframe/gpio_ie[15]
+ padframe/gpio_pullup[34] padframe/gpio_schmitt[35] padframe/gpio_out[3] padframe/gpio_out[0]
+ padframe/gpio_loopback_one[10] padframe/gpio_drive1[12] padframe/gpio_oe[5] padframe/gpio_slew[12]
+ padframe/gpio_slew[30] padframe/gpio_ie[37] padframe/gpio_ana[15] padframe/gpio_oe[2]
+ padframe/gpio_drive0[8] padframe/gpio_drive1[17] padframe/gpio_pullup[38] padframe/resetb_loopback_one
+ padframe/gpio_pulldown[12] padframe/gpio_drive1[34] padframe/gpio_pulldown[30] padframe/gpio_ie[16]
+ padframe/gpio_ie[34] padframe/gpio_loopback_one[33] padframe/gpio_slew[37] padframe/gpio_drive1[11]
+ padframe/mask_rev[27] gpio[0] padframe/gpio_pullup[17] padframe/mask_rev[29] padframe/gpio_in[20]
+ padframe/gpio_schmitt[18] padframe/gpio_pullup[35] padframe/gpio_schmitt[36] gpio[23]
+ padframe/gpio_out[8] padframe/gpio_ie[3] padframe/gpio_oe[9] padframe/gpio_slew[16]
+ padframe/gpio_ie[31] padframe/mask_rev[28] padframe/gpio_slew[34] padframe/gpio_out[5]
+ gpio[3] padframe/gpio_oe[37] padframe/gpio_slew[39] padframe/mask_rev[31] padframe/gpio_out[27]
+ padframe/gpio_drive0[38] padframe/gpio_out[2] padframe/gpio_out[24] padframe/gpio_in[40]
+ padframe/gpio_drive0[7] padframe/gpio_in[28] padframe/mask_rev[30] padframe/gpio_drive0[22]
+ padframe/gpio_in[22] padframe/gpio_drive1[16] gpio[42] padframe/gpio_oe[42] padframe/gpio_schmitt[33]
+ padframe/gpio_pulldown[19] gpio[20] padframe/gpio_pulldown[37] padframe/gpio_ie[0]
+ padframe/por_h padframe/gpio_oe[6] padframe/gpio_slew[13] padframe/gpio_ana[19]
+ padframe/gpio_slew[31] padframe/gpio_oe[25] padframe/gpio_oe[39] padframe/gpio_drive1[33]
+ gpio[41] padframe/gpio_loopback_zero[22] padframe/mask_rev[11] padframe/gpio_drive1[10]
+ padframe/gpio_ie[38] gpio[43] padframe/gpio_drive0[43] gpio[26] padframe/gpio_pulldown[6]
+ padframe/gpio_pullup[20] padframe/gpio_pullup[19] padframe/gpio_pullup[40] padframe/gpio_schmitt[21]
+ padframe/gpio_pulldown[16] padframe/gpio_out[21] padframe/gpio_pulldown[34] padframe/gpio_ie[41]
+ padframe/mask_rev[10] padframe/gpio_pulldown[39] padframe/gpio_drive0[27] padframe/mask_rev[13]
+ padframe/gpio_ana[16] padframe/gpio_oe[3] gpio[6] padframe/gpio_slew[10] padframe/gpio_oe[22]
+ padframe/gpio_schmitt[43] padframe/mask_rev[12] padframe/gpio_pullup[42] padframe/gpio_loopback_one[38]
+ padframe/mask_rev[15] padframe/gpio_schmitt[23] padframe/gpio_slew[38] padframe/gpio_drive0[6]
+ padframe/gpio_pulldown[3] padframe/gpio_pulldown[13] padframe/mask_rev[14] padframe/gpio_ie[7]
+ padframe/gpio_drive0[21] padframe/gpio_pulldown[31] padframe/gpio_ie[17] padframe/gpio_drive1[15]
+ padframe/gpio_ie[26] padframe/mask_rev[17] padframe/gpio_ie[35] padframe/gpio_drive1[39]
+ padframe/gpio_out[41] padframe/gpio_oe[0] padframe/gpio_drive1[0] padframe/mask_rev[16]
+ padframe/gpio_drive0[39] padframe/gpio_in[6] padframe/mask_rev[19] gpio[1] padframe/gpio_out[42]
+ padframe/gpio_drive1[32] padframe/gpio_slew[18] padframe/gpio_loopback_zero[41]
+ padframe/gpio_pullup[18] padframe/gpio_pullup[27] padframe/gpio_schmitt[19] padframe/gpio_pullup[36]
+ padframe/gpio_schmitt[28] padframe/gpio_schmitt[37] gpio[29] padframe/mask_rev[18]
+ padframe/gpio_oe[38] padframe/gpio_pulldown[0] padframe/gpio_pulldown[10] padframe/gpio_ie[4]
+ padframe/resetb_pullup padframe/gpio_ie[23] padframe/gpio_pullup[22] padframe/gpio_ie[32]
+ padframe/gpio_slew[17] padframe/gpio_oe[41] padframe/gpio_slew[35] padframe/gpio_oe[29]
+ gpio[9] padframe/gpio_pullup[39] gpio[14] padframe/gpio_out[43] padframe/gpio_out[7]
+ padframe/gpio_drive0[26] padframe/gpio_out[29] gpio[11] padframe/resetb_pulldown
+ padframe/gpio_schmitt[42] padframe/gpio_ana[20] padframe/gpio_out[4] padframe/gpio_pulldown[38]
+ padframe/gpio_out[26] padframe/gpio_loopback_zero[42] padframe/gpio_pullup[5] padframe/gpio_out[31]
+ padframe/gpio_drive1[5] padframe/gpio_pullup[24] padframe/gpio_ie[21] padframe/gpio_schmitt[16]
+ padframe/gpio_out[1] padframe/gpio_pulldown[41] gpio[24] padframe/gpio_schmitt[25]
+ gpio[40] padframe/gpio_schmitt[34] gpio[21] padframe/gpio_out[23] padframe/gpio_loopback_one[24]
+ padframe/gpio_loopback_zero[13] padframe/gpio_schmitt[39] padframe/gpio_drive1[20]
+ padframe/gpio_ie[1] padframe/gpio_drive1[37] padframe/gpio_out[15] padframe/gpio_ie[20]
+ padframe/gpio_ie[19] padframe/gpio_oe[7] padframe/gpio_slew[14] padframe/gpio_ie[40]
+ padframe/gpio_slew[23] padframe/gpio_out[20] gpio[4] padframe/gpio_slew[32] padframe/gpio_ana[39]
+ padframe/gpio_pulldown[20] padframe/gpio_oe[26] padframe/gpio_in[42] padframe/gpio_drive0[20]
+ padframe/gpio_drive1[14] padframe/gpio_out[12] gpio[31] padframe/gpio_drive0[37]
+ gpio[34] padframe/gpio_pulldown[18] padframe/gpio_loopback_one[42] gpio[8] padframe/gpio_pullup[2]
+ padframe/gpio_out[18] padframe/gpio_schmitt[3] padframe/gpio_ie[42] padframe/gpio_out[16]
+ padframe/gpio_pulldown[7] padframe/gpio_pullup[21] padframe/gpio_schmitt[22] padframe/gpio_pulldown[40]
+ padframe/gpio_slew[21] padframe/gpio_pulldown[17] padframe/gpio_schmitt[17] padframe/gpio_pulldown[26]
+ padframe/gpio_pulldown[35] padframe/gpio_drive1[31] padframe/gpio_slew[1] padframe/gpio_ana[17]
+ padframe/gpio_oe[4] padframe/gpio_slew[11] padframe/gpio_slew[20] padframe/gpio_slew[19]
+ padframe/gpio_slew[40] gpio[17] padframe/gpio_oe[14] vccd padframe/gpio_drive1[40]
+ padframe/gpio_in[23] padframe/gpio_oe[23] padframe/gpio_oe[32] padframe/gpio_in[21]
+ padframe/gpio_drive0[31] gpio[38] padframe/gpio_drive1[25] padframe/gpio_pullup[43]
+ gpio[18] padframe/gpio_loopback_one[39] padframe/gpio_pullup[23] padframe/gpio_drive0[40]
+ gpio[5] padframe/gpio_drive0[25] padframe/gpio_drive1[19] padframe/gpio_in[24] padframe/gpio_schmitt[41]
+ padframe/gpio_schmitt[0] gpio[27] padframe/gpio_pulldown[4] padframe/gpio_slew[42]
+ padframe/gpio_schmitt[10] padframe/gpio_pulldown[14] padframe/gpio_ie[8] padframe/gpio_pulldown[23]
+ gpio[28] padframe/gpio_pulldown[32] padframe/gpio_oe[21] padframe/gpio_ie[18] padframe/gpio_ie[27]
+ padframe/gpio_ie[36] padframe/gpio_ana[38] padframe/gpio_out[38] padframe/gpio_drive0[19]
+ padframe/gpio_drive1[4] gpio[7] padframe/gpio_oe[1] gpio[12] padframe/gpio_oe[11]
+ padframe/gpio_oe[20] padframe/gpio_oe[40] padframe/gpio_ie[22] padframe/gpio_drive1[36]
+ padframe/gpio_pullup[16] vddio padframe/gpio_ie[39] gpio[15] resetb padframe/gpio_drive0[4]
+ gpio[37] padframe/gpio_in[41] padframe/gpio_schmitt[38] padframe/gpio_out[40] vssd
+ gf180mcu_padframe
Xopenframe_project_wrapper_0 padframe/gpio_in[38] padframe/gpio_in[40] padframe/gpio_oe[40]
+ padframe/gpio_in[39] padframe/gpio_oe[39] padframe/gpio_in[41] padframe/gpio_out[41]
+ padframe/gpio_ie[41] padframe/gpio_oe[41] padframe/gpio_in[42] padframe/gpio_out[42]
+ padframe/gpio_ie[42] padframe/gpio_oe[42] padframe/gpio_drive0[38] padframe/gpio_drive2[38]
+ padframe/gpio_in[43] padframe/gpio_ie[38] padframe/gpio_out[38] padframe/gpio_oe[38]
+ padframe/gpio_pulldown[38] padframe/gpio_pullup[38] padframe/gpio_schmitt[38] padframe/gpio_slew[38]
+ padframe/gpio_schmitt[42] padframe/gpio_pullup[42] padframe/gpio_drive0[42] padframe/gpio_drive1[42]
+ padframe/gpio_pulldown[42] padframe/gpio_slew[42] padframe/gpio_schmitt[41] padframe/gpio_pullup[41]
+ padframe/gpio_drive0[41] padframe/gpio_drive1[41] padframe/gpio_pulldown[41] padframe/gpio_slew[41]
+ padframe/gpio_schmitt[40] padframe/gpio_pullup[40] padframe/gpio_drive0[40] padframe/gpio_drive1[40]
+ padframe/gpio_pulldown[40] padframe/gpio_ie[40] padframe/gpio_slew[40] padframe/gpio_out[40]
+ padframe/gpio_schmitt[39] padframe/gpio_pullup[39] padframe/gpio_drive0[39] padframe/gpio_drive1[39]
+ padframe/gpio_pulldown[39] padframe/gpio_ie[39] padframe/gpio_slew[39] padframe/gpio_out[39]
+ padframe/gpio_out[43] padframe/gpio_slew[43] padframe/gpio_ie[43] padframe/gpio_pulldown[43]
+ padframe/gpio_drive1[43] padframe/gpio_drive0[43] padframe/gpio_pullup[43] padframe/gpio_schmitt[43]
+ padframe/gpio_oe[43] padframe/gpio_drive0[30] padframe/gpio_drive0[0] padframe/gpio_drive0[5]
+ padframe/gpio_drive1[5] padframe/gpio_drive0[6] padframe/gpio_drive1[6] padframe/gpio_drive0[7]
+ padframe/gpio_drive1[7] padframe/gpio_drive0[8] padframe/gpio_drive1[8] padframe/gpio_drive0[9]
+ padframe/gpio_drive1[9] padframe/gpio_drive1[0] padframe/gpio_drive0[10] padframe/gpio_drive1[10]
+ padframe/gpio_drive0[11] padframe/gpio_drive1[11] padframe/gpio_drive0[12] padframe/gpio_drive1[12]
+ padframe/gpio_drive0[13] padframe/gpio_drive1[13] padframe/gpio_drive0[14] padframe/gpio_drive1[14]
+ padframe/gpio_drive0[1] padframe/gpio_drive0[15] padframe/gpio_drive1[15] padframe/gpio_drive0[16]
+ padframe/gpio_drive1[16] padframe/gpio_drive0[17] padframe/gpio_drive1[17] padframe/gpio_drive0[18]
+ padframe/gpio_drive1[18] padframe/gpio_drive0[19] padframe/gpio_drive1[1] padframe/gpio_drive0[20]
+ padframe/gpio_drive1[20] padframe/gpio_drive0[21] padframe/gpio_drive1[21] padframe/gpio_drive0[22]
+ padframe/gpio_drive1[22] padframe/gpio_drive0[23] padframe/gpio_drive1[23] padframe/gpio_drive0[24]
+ padframe/gpio_drive1[24] padframe/gpio_drive0[2] padframe/gpio_drive1[25] padframe/gpio_drive0[25]
+ padframe/gpio_drive0[26] padframe/gpio_drive1[26] padframe/gpio_drive0[27] padframe/gpio_drive1[27]
+ padframe/gpio_drive0[28] padframe/gpio_drive1[28] padframe/gpio_drive0[29] padframe/gpio_drive1[29]
+ padframe/gpio_drive1[2] padframe/gpio_drive1[30] padframe/gpio_drive0[31] padframe/gpio_drive1[31]
+ padframe/gpio_drive0[32] padframe/gpio_drive1[32] padframe/gpio_drive0[33] padframe/gpio_drive1[33]
+ padframe/gpio_drive0[34] padframe/gpio_drive1[34] padframe/gpio_drive0[3] padframe/gpio_drive0[35]
+ padframe/gpio_drive1[35] padframe/gpio_drive0[36] padframe/gpio_drive1[36] padframe/gpio_drive0[37]
+ padframe/gpio_drive1[37] padframe/gpio_drive1[3] padframe/gpio_drive0[4] padframe/gpio_drive1[4]
+ padframe/gpio_in[0] padframe/gpio_in[10] padframe/gpio_in[11] padframe/gpio_in[12]
+ padframe/gpio_in[13] padframe/gpio_in[14] padframe/gpio_in[15] padframe/gpio_in[16]
+ padframe/gpio_in[17] padframe/gpio_in[18] padframe/gpio_in[19] padframe/gpio_in[1]
+ padframe/gpio_in[20] padframe/gpio_in[21] padframe/gpio_in[22] padframe/gpio_in[23]
+ padframe/gpio_in[24] padframe/gpio_in[25] padframe/gpio_in[26] padframe/gpio_in[27]
+ padframe/gpio_in[28] padframe/gpio_in[29] padframe/gpio_in[2] padframe/gpio_in[30]
+ padframe/gpio_in[31] padframe/gpio_in[32] padframe/gpio_in[33] padframe/gpio_in[34]
+ padframe/gpio_in[35] padframe/gpio_in[36] padframe/gpio_in[37] padframe/gpio_in[3]
+ padframe/gpio_in[4] padframe/gpio_in[5] padframe/gpio_in[6] padframe/gpio_in[7]
+ padframe/gpio_in[8] padframe/gpio_in[9] padframe/gpio_ie[0] padframe/gpio_ie[10]
+ padframe/gpio_ie[11] padframe/gpio_ie[12] padframe/gpio_ie[13] padframe/gpio_ie[14]
+ padframe/gpio_ie[15] padframe/gpio_ie[16] padframe/gpio_ie[17] padframe/gpio_ie[18]
+ padframe/gpio_ie[19] padframe/gpio_ie[1] padframe/gpio_ie[20] padframe/gpio_ie[21]
+ padframe/gpio_ie[22] padframe/gpio_ie[23] padframe/gpio_ie[24] padframe/gpio_ie[25]
+ padframe/gpio_ie[26] padframe/gpio_ie[27] padframe/gpio_ie[28] padframe/gpio_ie[29]
+ padframe/gpio_ie[2] padframe/gpio_ie[30] padframe/gpio_ie[31] padframe/gpio_ie[32]
+ padframe/gpio_ie[33] padframe/gpio_ie[34] padframe/gpio_ie[35] padframe/gpio_ie[36]
+ padframe/gpio_ie[37] padframe/gpio_ie[3] padframe/gpio_ie[4] padframe/gpio_ie[5]
+ padframe/gpio_ie[6] padframe/gpio_ie[7] padframe/gpio_ie[8] padframe/gpio_ie[9]
+ padframe/gpio_out[0] padframe/gpio_out[10] padframe/gpio_out[11] padframe/gpio_out[12]
+ padframe/gpio_out[13] padframe/gpio_out[14] padframe/gpio_out[15] padframe/gpio_out[16]
+ padframe/gpio_out[17] padframe/gpio_out[18] padframe/gpio_out[19] padframe/gpio_out[1]
+ padframe/gpio_out[20] padframe/gpio_out[21] padframe/gpio_out[22] padframe/gpio_out[23]
+ padframe/gpio_out[24] padframe/gpio_out[25] padframe/gpio_out[26] padframe/gpio_out[27]
+ padframe/gpio_out[28] padframe/gpio_out[29] padframe/gpio_out[2] padframe/gpio_out[30]
+ padframe/gpio_out[31] padframe/gpio_out[32] padframe/gpio_out[33] padframe/gpio_out[34]
+ padframe/gpio_out[35] padframe/gpio_out[36] padframe/gpio_out[37] padframe/gpio_out[3]
+ padframe/gpio_out[4] padframe/gpio_out[5] padframe/gpio_out[6] padframe/gpio_out[7]
+ padframe/gpio_out[8] padframe/gpio_out[9] padframe/gpio_oe[0] padframe/gpio_oe[10]
+ padframe/gpio_oe[11] padframe/gpio_oe[12] padframe/gpio_oe[13] padframe/gpio_oe[14]
+ padframe/gpio_oe[15] padframe/gpio_oe[16] padframe/gpio_oe[17] padframe/gpio_oe[18]
+ padframe/gpio_oe[19] padframe/gpio_oe[1] padframe/gpio_oe[20] padframe/gpio_oe[21]
+ padframe/gpio_oe[22] padframe/gpio_oe[23] padframe/gpio_oe[24] padframe/gpio_oe[25]
+ padframe/gpio_oe[26] padframe/gpio_oe[27] padframe/gpio_oe[28] padframe/gpio_oe[29]
+ padframe/gpio_oe[2] padframe/gpio_oe[30] padframe/gpio_oe[31] padframe/gpio_oe[32]
+ padframe/gpio_oe[33] padframe/gpio_oe[34] padframe/gpio_oe[35] padframe/gpio_oe[36]
+ padframe/gpio_oe[37] padframe/gpio_oe[3] padframe/gpio_oe[4] padframe/gpio_oe[5]
+ padframe/gpio_oe[6] padframe/gpio_oe[7] padframe/gpio_oe[8] padframe/gpio_oe[9]
+ padframe/gpio_pulldown[0] padframe/gpio_pulldown[10] padframe/gpio_pulldown[11]
+ padframe/gpio_pulldown[12] padframe/gpio_pulldown[13] padframe/gpio_pulldown[14]
+ padframe/gpio_pulldown[15] padframe/gpio_pulldown[16] padframe/gpio_pulldown[17]
+ padframe/gpio_pulldown[18] padframe/gpio_pulldown[19] padframe/gpio_pulldown[1]
+ padframe/gpio_pulldown[20] padframe/gpio_pulldown[21] padframe/gpio_pulldown[22]
+ padframe/gpio_pulldown[23] padframe/gpio_pulldown[24] padframe/gpio_pulldown[25]
+ padframe/gpio_pulldown[26] padframe/gpio_pulldown[27] padframe/gpio_pulldown[28]
+ padframe/gpio_pulldown[29] padframe/gpio_pulldown[2] padframe/gpio_pulldown[30]
+ padframe/gpio_pulldown[31] padframe/gpio_pulldown[32] padframe/gpio_pulldown[33]
+ padframe/gpio_pulldown[34] padframe/gpio_pulldown[35] padframe/gpio_pulldown[36]
+ padframe/gpio_pulldown[37] padframe/gpio_pulldown[3] padframe/gpio_pulldown[4] padframe/gpio_pulldown[5]
+ padframe/gpio_pulldown[6] padframe/gpio_pulldown[7] padframe/gpio_pulldown[8] padframe/gpio_pulldown[9]
+ padframe/gpio_pullup[0] padframe/gpio_pullup[10] padframe/gpio_pullup[11] padframe/gpio_pullup[12]
+ padframe/gpio_pullup[13] padframe/gpio_pullup[14] padframe/gpio_pullup[15] padframe/gpio_pullup[16]
+ padframe/gpio_pullup[17] padframe/gpio_pullup[18] padframe/gpio_pullup[19] padframe/gpio_pullup[1]
+ padframe/gpio_pullup[20] padframe/gpio_pullup[21] padframe/gpio_pullup[22] padframe/gpio_pullup[23]
+ padframe/gpio_pullup[24] padframe/gpio_pullup[25] padframe/gpio_pullup[26] padframe/gpio_pullup[27]
+ padframe/gpio_pullup[28] padframe/gpio_pullup[29] padframe/gpio_pullup[2] padframe/gpio_pullup[30]
+ padframe/gpio_pullup[31] padframe/gpio_pullup[32] padframe/gpio_pullup[33] padframe/gpio_pullup[34]
+ padframe/gpio_pullup[35] padframe/gpio_pullup[36] padframe/gpio_pullup[37] padframe/gpio_pullup[3]
+ padframe/gpio_pullup[4] padframe/gpio_pullup[5] padframe/gpio_pullup[6] padframe/gpio_pullup[7]
+ padframe/gpio_pullup[8] padframe/gpio_pullup[9] padframe/gpio_schmitt[0] padframe/gpio_schmitt[10]
+ padframe/gpio_schmitt[11] padframe/gpio_schmitt[12] padframe/gpio_schmitt[13] padframe/gpio_schmitt[14]
+ padframe/gpio_schmitt[15] padframe/gpio_schmitt[16] padframe/gpio_schmitt[17] padframe/gpio_schmitt[18]
+ padframe/gpio_schmitt[19] padframe/gpio_schmitt[1] padframe/gpio_schmitt[20] padframe/gpio_schmitt[21]
+ padframe/gpio_schmitt[22] padframe/gpio_schmitt[23] padframe/gpio_schmitt[24] padframe/gpio_schmitt[25]
+ padframe/gpio_schmitt[26] padframe/gpio_schmitt[27] padframe/gpio_schmitt[28] padframe/gpio_schmitt[29]
+ padframe/gpio_schmitt[2] padframe/gpio_schmitt[30] padframe/gpio_schmitt[31] padframe/gpio_schmitt[32]
+ padframe/gpio_schmitt[33] padframe/gpio_schmitt[34] padframe/gpio_schmitt[35] padframe/gpio_schmitt[36]
+ padframe/gpio_schmitt[37] padframe/gpio_schmitt[3] padframe/gpio_schmitt[4] padframe/gpio_schmitt[5]
+ padframe/gpio_schmitt[6] padframe/gpio_schmitt[7] padframe/gpio_schmitt[8] padframe/gpio_schmitt[9]
+ padframe/gpio_slew[0] padframe/gpio_slew[10] padframe/gpio_slew[11] padframe/gpio_slew[12]
+ padframe/gpio_slew[13] padframe/gpio_slew[14] padframe/gpio_slew[15] padframe/gpio_slew[16]
+ padframe/gpio_slew[17] padframe/gpio_slew[18] padframe/gpio_slew[19] padframe/gpio_slew[1]
+ padframe/gpio_slew[20] padframe/gpio_slew[21] padframe/gpio_slew[22] padframe/gpio_slew[23]
+ padframe/gpio_slew[24] padframe/gpio_slew[25] padframe/gpio_slew[26] padframe/gpio_slew[27]
+ padframe/gpio_slew[28] padframe/gpio_slew[29] padframe/gpio_slew[2] padframe/gpio_slew[30]
+ padframe/gpio_slew[31] padframe/gpio_slew[32] padframe/gpio_slew[33] padframe/gpio_slew[34]
+ padframe/gpio_slew[35] padframe/gpio_slew[36] padframe/gpio_slew[37] padframe/gpio_slew[3]
+ padframe/gpio_slew[4] padframe/gpio_slew[5] padframe/gpio_slew[6] padframe/gpio_slew[7]
+ padframe/gpio_slew[8] padframe/gpio_slew[9] padframe/resetb_core padframe/gpio_ana[0]
+ padframe/gpio_ana[1] padframe/gpio_ana[2] padframe/gpio_ana[3] padframe/gpio_ana[4]
+ padframe/gpio_ana[5] padframe/gpio_ana[6] padframe/gpio_ana[7] padframe/gpio_ana[8]
+ padframe/gpio_ana[9] padframe/gpio_ana[10] padframe/gpio_ana[11] padframe/gpio_ana[12]
+ padframe/gpio_ana[13] padframe/gpio_ana[14] padframe/gpio_ana[15] padframe/gpio_ana[16]
+ padframe/gpio_ana[17] padframe/gpio_ana[18] padframe/gpio_ana[19] padframe/gpio_ana[20]
+ padframe/gpio_ana[21] padframe/gpio_ana[22] padframe/gpio_ana[23] padframe/gpio_ana[24]
+ padframe/gpio_ana[25] padframe/gpio_ana[26] padframe/gpio_ana[27] padframe/gpio_ana[28]
+ padframe/gpio_ana[29] padframe/gpio_ana[30] padframe/gpio_ana[31] padframe/gpio_ana[32]
+ padframe/gpio_ana[33] padframe/gpio_ana[34] padframe/gpio_ana[35] padframe/gpio_ana[36]
+ padframe/gpio_ana[37] padframe/gpio_ana[38] padframe/gpio_ana[39] padframe/gpio_ana[40]
+ padframe/gpio_ana[41] padframe/gpio_ana[42] padframe/gpio_ana[43] padframe/gpio_loopback_zero[0]
+ padframe/gpio_loopback_one[0] padframe/gpio_loopback_zero[1] padframe/gpio_loopback_one[1]
+ padframe/gpio_loopback_zero[2] padframe/gpio_loopback_one[2] padframe/gpio_loopback_one[3]
+ padframe/gpio_loopback_zero[3] padframe/gpio_loopback_zero[4] padframe/gpio_loopback_one[4]
+ padframe/gpio_loopback_one[5] padframe/gpio_loopback_zero[5] padframe/gpio_loopback_zero[6]
+ padframe/gpio_loopback_one[6] padframe/gpio_loopback_one[7] padframe/gpio_loopback_zero[7]
+ padframe/gpio_loopback_zero[8] padframe/gpio_loopback_one[8] padframe/gpio_loopback_one[9]
+ padframe/gpio_loopback_zero[9] padframe/gpio_loopback_zero[10] padframe/gpio_loopback_one[10]
+ padframe/gpio_loopback_one[11] padframe/gpio_loopback_zero[11] padframe/gpio_loopback_zero[12]
+ padframe/gpio_loopback_one[12] padframe/gpio_loopback_one[13] padframe/gpio_loopback_zero[14]
+ padframe/gpio_loopback_one[14] padframe/gpio_loopback_one[15] padframe/gpio_loopback_zero[15]
+ padframe/gpio_loopback_zero[16] padframe/gpio_loopback_one[16] padframe/gpio_loopback_one[17]
+ padframe/gpio_loopback_zero[17] padframe/gpio_loopback_zero[18] padframe/gpio_loopback_one[18]
+ padframe/gpio_loopback_one[19] padframe/gpio_loopback_zero[19] padframe/gpio_loopback_zero[20]
+ padframe/gpio_loopback_one[20] padframe/gpio_loopback_one[21] padframe/gpio_loopback_zero[21]
+ padframe/gpio_loopback_zero[22] padframe/gpio_loopback_one[22] padframe/gpio_loopback_one[23]
+ padframe/gpio_loopback_zero[23] padframe/gpio_loopback_zero[24] padframe/gpio_loopback_one[24]
+ padframe/gpio_loopback_one[25] padframe/gpio_loopback_zero[25] padframe/gpio_loopback_zero[26]
+ padframe/gpio_loopback_one[26] padframe/gpio_loopback_one[27] padframe/gpio_loopback_zero[27]
+ padframe/gpio_loopback_zero[28] padframe/gpio_loopback_one[28] padframe/gpio_loopback_one[29]
+ padframe/gpio_loopback_zero[29] padframe/gpio_loopback_zero[30] padframe/gpio_loopback_one[30]
+ padframe/gpio_loopback_one[31] padframe/gpio_loopback_zero[31] padframe/gpio_loopback_zero[32]
+ padframe/gpio_loopback_one[32] padframe/gpio_loopback_one[33] padframe/gpio_loopback_zero[33]
+ padframe/gpio_loopback_zero[34] padframe/gpio_loopback_one[34] padframe/gpio_loopback_one[35]
+ padframe/gpio_loopback_zero[35] padframe/gpio_loopback_zero[36] padframe/gpio_loopback_one[36]
+ padframe/gpio_loopback_one[37] padframe/gpio_loopback_zero[37] padframe/gpio_loopback_zero[38]
+ padframe/gpio_loopback_one[38] padframe/gpio_loopback_one[39] padframe/gpio_loopback_zero[39]
+ padframe/gpio_loopback_zero[40] padframe/gpio_loopback_one[40] padframe/gpio_loopback_one[41]
+ padframe/gpio_loopback_zero[41] padframe/gpio_loopback_zero[42] padframe/gpio_loopback_one[42]
+ padframe/gpio_loopback_one[43] padframe/gpio_loopback_zero[43] padframe/resetb_pullup
+ padframe/resetb_pulldown padframe/resetb_loopback_one padframe/resetb_loopback_zero
+ padframe/por_h padframe/porb_h padframe/porb_l padframe/mask_rev[0] padframe/mask_rev[1]
+ padframe/mask_rev[2] padframe/mask_rev[3] padframe/mask_rev[4] padframe/mask_rev[5]
+ padframe/mask_rev[6] padframe/mask_rev[7] padframe/mask_rev[8] padframe/mask_rev[9]
+ padframe/mask_rev[10] padframe/mask_rev[11] padframe/mask_rev[12] padframe/mask_rev[13]
+ padframe/mask_rev[14] padframe/mask_rev[15] padframe/mask_rev[16] padframe/mask_rev[17]
+ padframe/mask_rev[18] padframe/mask_rev[19] padframe/mask_rev[20] padframe/mask_rev[21]
+ padframe/mask_rev[22] padframe/mask_rev[23] padframe/mask_rev[24] padframe/mask_rev[25]
+ padframe/mask_rev[26] padframe/mask_rev[27] padframe/mask_rev[28] padframe/mask_rev[29]
+ padframe/mask_rev[30] padframe/mask_rev[31] vssd vssd vddio vccd padframe/gpio_pulldown[7]
+ padframe/gpio_schmitt[5] padframe/gpio_pulldown[5] padframe/gpio_ie[10] padframe/gpio_slew[25]
+ padframe/gpio_slew[28] padframe/gpio_schmitt[0] padframe/gpio_pulldown[0] padframe/gpio_ie[3]
+ padframe/gpio_slew[24] padframe/gpio_slew[27] padframe/gpio_drive0[29] padframe/gpio_drive1[12]
+ padframe/gpio_ie[25] padframe/gpio_drive0[34] padframe/gpio_slew[0] padframe/gpio_drive1[7]
+ padframe/gpio_drive1[5] padframe/gpio_pullup[11] padframe/gpio_slew[1] padframe/gpio_drive1[0]
+ padframe/gpio_pulldown[29] padframe/gpio_schmitt[29] padframe/gpio_pullup[4] padframe/gpio_schmitt[34]
+ padframe/gpio_pulldown[34] padframe/gpio_slew[2] padframe/gpio_pullup[24] padframe/gpio_ie[31]
+ padframe/gpio_slew[3] padframe/gpio_ie[37] padframe/gpio_drive0[11] padframe/gpio_drive1[29]
+ padframe/gpio_slew[4] padframe/gpio_drive0[4] padframe/gpio_drive1[34] padframe/gpio_pullup[30]
+ padframe/gpio_slew[5] padframe/gpio_drive0[24] padframe/gpio_pullup[36] padframe/gpio_schmitt[11]
+ padframe/gpio_pulldown[11] padframe/gpio_slew[6] padframe/gpio_ie[14] padframe/gpio_pulldown[4]
+ padframe/gpio_schmitt[4] padframe/gpio_ie[9] padframe/gpio_schmitt[24] padframe/gpio_pulldown[24]
+ padframe/gpio_ie[2] padframe/gpio_drive0[30] padframe/gpio_drive1[11] padframe/gpio_pullup[35]
+ padframe/gpio_ie[26] padframe/gpio_drive0[36] padframe/gpio_drive1[4] padframe/gpio_pullup[10]
+ padframe/gpio_drive1[24] padframe/gpio_schmitt[30] padframe/gpio_pulldown[30] padframe/gpio_pullup[3]
+ padframe/gpio_ie[27] padframe/gpio_schmitt[36] padframe/gpio_pulldown[36] padframe/gpio_pullup[25]
+ padframe/gpio_ie[32] padframe/gpio_drive0[35] padframe/gpio_drive0[10] padframe/gpio_drive1[30]
+ padframe/gpio_drive0[3] padframe/gpio_drive1[36] padframe/gpio_pullup[31] padframe/gpio_schmitt[35]
+ padframe/gpio_pulldown[35] padframe/gpio_drive0[25] padframe/gpio_pullup[37] padframe/gpio_schmitt[10]
+ padframe/gpio_pulldown[10] padframe/gpio_ie[13] padframe/gpio_pulldown[3] padframe/gpio_schmitt[3]
+ padframe/gpio_ie[8] padframe/gpio_ie[6] padframe/gpio_schmitt[25] padframe/gpio_pulldown[25]
+ padframe/gpio_drive1[19] padframe/gpio_drive1[35] padframe/gpio_ie[1] padframe/gpio_drive0[31]
+ padframe/gpio_drive1[10] padframe/gpio_pullup[14] padframe/gpio_drive0[37] padframe/gpio_drive1[3]
+ padframe/gpio_pullup[9] padframe/gpio_drive1[25] padframe/gpio_schmitt[31] padframe/gpio_pullup[2]
+ padframe/gpio_pulldown[31] padframe/gpio_ie[28] padframe/gpio_schmitt[37] padframe/gpio_pulldown[37]
+ padframe/gpio_pullup[26] padframe/gpio_ie[33] padframe/gpio_drive0[14] padframe/gpio_drive0[9]
+ padframe/gpio_drive1[31] padframe/gpio_pullup[27] padframe/gpio_drive0[2] padframe/gpio_drive1[37]
+ padframe/gpio_pullup[32] padframe/gpio_schmitt[14] padframe/gpio_pulldown[14] padframe/gpio_drive0[26]
+ padframe/gpio_oe[7] padframe/gpio_schmitt[9] padframe/gpio_pulldown[9] padframe/gpio_out[7]
+ padframe/gpio_ie[12] padframe/gpio_schmitt[2] padframe/gpio_oe[8] padframe/gpio_pulldown[2]
+ padframe/gpio_out[8] padframe/gpio_ie[7] padframe/gpio_ie[5] padframe/gpio_drive0[27]
+ padframe/gpio_schmitt[26] padframe/gpio_pulldown[26] padframe/gpio_drive1[14] padframe/gpio_oe[9]
+ padframe/gpio_oe[37] padframe/gpio_out[9] padframe/gpio_out[37] padframe/gpio_ie[0]
+ padframe/gpio_drive0[32] padframe/gpio_drive1[9] padframe/gpio_oe[10] padframe/gpio_pullup[13]
+ padframe/gpio_oe[36] padframe/gpio_out[10] padframe/gpio_out[36] padframe/gpio_drive1[2]
+ padframe/gpio_pullup[8] padframe/gpio_schmitt[27] padframe/gpio_pullup[6] padframe/gpio_pulldown[27]
+ padframe/gpio_oe[11] padframe/gpio_oe[34] padframe/gpio_out[11] padframe/gpio_out[34]
+ padframe/gpio_drive1[26] padframe/gpio_schmitt[32] padframe/gpio_pulldown[32] padframe/gpio_pullup[1]
+ padframe/gpio_oe[12] padframe/gpio_ie[29] padframe/gpio_oe[33] padframe/gpio_out[12]
+ padframe/gpio_out[33] padframe/gpio_ie[34] padframe/gpio_oe[13] padframe/gpio_out[13]
+ padframe/gpio_oe[32] padframe/gpio_out[32] padframe/gpio_drive0[13] padframe/gpio_drive1[27]
+ padframe/gpio_oe[14] padframe/gpio_drive0[8] padframe/gpio_drive0[6] padframe/gpio_oe[31]
+ padframe/gpio_out[14] padframe/gpio_drive1[32] padframe/gpio_out[31] padframe/gpio_pullup[28]
+ padframe/gpio_drive0[1] padframe/gpio_oe[35] padframe/gpio_oe[30] padframe/gpio_out[35]
+ padframe/gpio_pullup[33] padframe/gpio_out[30] padframe/gpio_schmitt[13] padframe/gpio_pulldown[13]
+ padframe/gpio_slew[7] padframe/gpio_oe[26] padframe/gpio_schmitt[8] padframe/gpio_oe[29]
+ padframe/gpio_pulldown[8] padframe/gpio_out[26] padframe/gpio_out[29] padframe/gpio_schmitt[6]
+ padframe/gpio_pulldown[6] padframe/gpio_ie[11] padframe/gpio_slew[8] padframe/gpio_oe[25]
+ padframe/gpio_schmitt[1] padframe/gpio_oe[28] padframe/gpio_pulldown[1] padframe/gpio_out[25]
+ padframe/gpio_out[28] padframe/gpio_ie[4] padframe/gpio_slew[9] padframe/gpio_drive0[28]
+ padframe/gpio_slew[37] padframe/gpio_oe[27] padframe/gpio_drive1[13] padframe/gpio_oe[24]
+ padframe/gpio_out[24] padframe/gpio_out[27] padframe/gpio_ie[24] padframe/gpio_drive0[33]
+ padframe/gpio_slew[10] padframe/gpio_slew[36] padframe/gpio_drive1[8] padframe/gpio_drive1[6]
+ padframe/gpio_oe[0] padframe/gpio_pullup[12] padframe/gpio_out[0] padframe/gpio_slew[11]
+ padframe/gpio_drive1[1] padframe/gpio_pullup[7] padframe/gpio_slew[34] padframe/gpio_schmitt[28]
+ padframe/gpio_pulldown[28] padframe/gpio_pullup[5] padframe/gpio_oe[1] padframe/gpio_out[1]
+ padframe/gpio_schmitt[33] padframe/gpio_slew[12] padframe/gpio_pulldown[33] padframe/gpio_slew[33]
+ padframe/gpio_loopback_zero[13] padframe/gpio_pullup[0] padframe/gpio_oe[2] padframe/gpio_out[2]
+ padframe/gpio_ie[30] padframe/gpio_slew[13] padframe/gpio_slew[32] padframe/gpio_ie[36]
+ padframe/gpio_oe[3] padframe/gpio_out[3] padframe/gpio_drive0[12] padframe/gpio_drive1[28]
+ padframe/gpio_slew[14] padframe/gpio_slew[31] padframe/gpio_oe[4] padframe/gpio_drive0[7]
+ padframe/gpio_out[4] padframe/gpio_drive0[5] padframe/gpio_drive1[33] padframe/gpio_pullup[29]
+ padframe/gpio_slew[35] padframe/gpio_slew[30] padframe/gpio_drive0[0] padframe/gpio_oe[5]
+ padframe/gpio_out[5] padframe/gpio_pullup[34] padframe/gpio_schmitt[12] padframe/gpio_pulldown[12]
+ padframe/gpio_slew[26] padframe/gpio_slew[29] padframe/gpio_ie[35] padframe/gpio_oe[6]
+ padframe/gpio_schmitt[7] padframe/gpio_out[6] openframe_project_wrapper
.ends

