magic
tech gf180mcuD
magscale 1 5
timestamp 1766953626
<< metal1 >>
rect 0 489 30 519
<< via1 >>
rect 194 489 224 519
rect 866 489 896 519
rect 1426 489 1456 519
rect 2098 489 2128 519
rect 2658 489 2688 519
rect 3330 489 3360 519
rect 3890 489 3920 519
rect 4562 489 4592 519
rect 5122 489 5152 519
rect 5794 489 5824 519
rect 6354 489 6384 519
rect 7026 489 7056 519
rect 7586 489 7616 519
rect 8258 489 8288 519
rect 8818 489 8848 519
rect 9490 489 9520 519
rect 194 0 224 30
rect 866 0 896 30
rect 1426 0 1456 30
rect 2098 0 2128 30
rect 2658 0 2688 30
rect 3330 0 3360 30
rect 3890 0 3920 30
rect 4562 0 4592 30
rect 5122 0 5152 30
rect 5794 0 5824 30
rect 6354 0 6384 30
rect 7026 0 7056 30
rect 7586 0 7616 30
rect 8258 0 8288 30
rect 8818 0 8848 30
rect 9490 0 9520 30
<< properties >>
string flatten true
<< end >>
