VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ring_osc2x13
  CLASS BLOCK ;
  FOREIGN ring_osc2x13 ;
  ORIGIN 6.810 -16.710 ;
  SIZE 68.060 BY 56.035 ;
  PIN vdd
    ANTENNADIFFAREA 382.877380 ;
    PORT
      LAYER Nwell ;
        RECT -6.810 71.745 60.970 72.450 ;
        RECT -6.810 69.870 -5.810 71.745 ;
        RECT 60.250 69.870 60.970 71.745 ;
        RECT -6.810 62.030 -5.810 66.330 ;
        RECT 60.250 62.030 61.250 66.330 ;
        RECT -6.810 54.190 -5.810 58.490 ;
        RECT 60.250 54.190 61.250 58.490 ;
        RECT -6.810 46.350 -5.810 50.650 ;
        RECT 60.250 46.350 61.250 50.650 ;
        RECT -6.810 38.510 -5.810 42.810 ;
        RECT 60.250 38.510 61.250 42.810 ;
        RECT -6.810 30.670 -5.810 34.970 ;
        RECT 60.250 30.670 61.250 34.970 ;
        RECT -6.810 22.830 -5.810 27.130 ;
        RECT 60.250 22.830 61.250 27.130 ;
        RECT -6.810 17.710 -5.810 19.290 ;
        RECT 60.250 17.710 61.250 19.290 ;
        RECT -6.810 16.710 61.250 17.710 ;
      LAYER Metal1 ;
        RECT -6.380 71.745 60.540 72.320 ;
        RECT -6.380 71.720 -5.810 71.745 ;
        RECT 60.250 71.720 60.540 71.745 ;
        RECT -6.005 70.335 -5.810 71.720 ;
        RECT -5.975 64.480 -5.810 65.865 ;
        RECT 60.250 64.480 60.445 65.865 ;
        RECT -6.380 63.880 -1.900 64.480 ;
        RECT 60.250 63.880 60.820 64.480 ;
        RECT -6.005 62.495 -5.810 63.880 ;
        RECT 60.250 62.495 60.415 63.880 ;
        RECT -6.005 56.640 -5.810 58.025 ;
        RECT -6.380 56.040 -5.810 56.640 ;
        RECT -5.975 54.655 -5.810 56.040 ;
        RECT 60.250 56.640 60.415 58.025 ;
        RECT 60.250 56.040 60.820 56.640 ;
        RECT 60.250 54.655 60.445 56.040 ;
        RECT -5.975 48.800 -5.810 50.185 ;
        RECT -6.380 48.200 -5.810 48.800 ;
        RECT -6.005 46.815 -5.810 48.200 ;
        RECT 60.250 48.800 60.445 50.185 ;
        RECT 60.250 48.200 60.820 48.800 ;
        RECT 60.250 46.815 60.415 48.200 ;
        RECT -6.005 40.960 -5.810 42.345 ;
        RECT -6.380 40.360 -5.810 40.960 ;
        RECT -5.975 38.975 -5.810 40.360 ;
        RECT 60.250 40.960 60.415 42.345 ;
        RECT 60.250 40.360 60.820 40.960 ;
        RECT 60.250 38.975 60.445 40.360 ;
        RECT -5.975 33.120 -5.810 34.505 ;
        RECT -6.380 32.520 -5.810 33.120 ;
        RECT -6.005 31.135 -5.810 32.520 ;
        RECT 60.250 33.120 60.445 34.505 ;
        RECT 60.250 32.520 60.820 33.120 ;
        RECT 60.250 31.135 60.415 32.520 ;
        RECT -6.005 25.280 -5.810 26.665 ;
        RECT -6.380 24.680 -5.810 25.280 ;
        RECT -5.975 23.295 -5.810 24.680 ;
        RECT 60.250 25.280 60.415 26.665 ;
        RECT 60.250 24.680 60.820 25.280 ;
        RECT 60.250 23.295 60.445 24.680 ;
        RECT -6.005 17.710 -5.810 18.825 ;
        RECT 60.250 17.710 60.415 18.825 ;
        RECT -6.005 17.440 -5.665 17.710 ;
        RECT -3.935 17.440 -3.705 17.710 ;
        RECT -1.695 17.440 -1.465 17.710 ;
        RECT 1.475 17.440 1.705 17.710 ;
        RECT 3.925 17.440 4.155 17.710 ;
        RECT 7.965 17.440 8.195 17.710 ;
        RECT 10.435 17.440 10.665 17.710 ;
        RECT 12.885 17.440 13.115 17.710 ;
        RECT 16.925 17.440 17.155 17.710 ;
        RECT 18.465 17.440 18.695 17.710 ;
        RECT 20.065 17.440 20.295 17.710 ;
        RECT 21.635 17.440 21.865 17.710 ;
        RECT 24.085 17.440 24.315 17.710 ;
        RECT 28.125 17.440 28.355 17.710 ;
        RECT 29.865 17.440 30.205 17.710 ;
        RECT 31.715 17.440 31.945 17.710 ;
        RECT 34.165 17.440 34.395 17.710 ;
        RECT 38.205 17.440 38.435 17.710 ;
        RECT 40.145 17.440 40.375 17.710 ;
        RECT 41.745 17.440 41.975 17.710 ;
        RECT 43.345 17.440 43.575 17.710 ;
        RECT 45.185 17.440 45.415 17.710 ;
        RECT 46.785 17.440 47.015 17.710 ;
        RECT 48.385 17.440 48.615 17.710 ;
        RECT 49.825 17.440 50.055 17.710 ;
        RECT 51.425 17.440 51.655 17.710 ;
        RECT 52.065 17.440 52.295 17.710 ;
        RECT 53.665 17.440 53.895 17.710 ;
        RECT 54.305 17.440 54.535 17.710 ;
        RECT 56.545 17.440 56.775 17.710 ;
        RECT 60.075 17.440 60.415 17.710 ;
        RECT -6.380 16.840 60.820 17.440 ;
      LAYER Metal2 ;
        RECT -0.835 71.745 0.250 72.330 ;
        RECT 23.895 71.745 24.960 72.330 ;
        RECT 38.370 71.745 39.430 72.335 ;
        RECT -0.790 17.440 0.200 17.710 ;
        RECT 24.190 17.440 25.180 17.710 ;
        RECT 39.095 17.440 40.085 17.710 ;
        RECT -0.835 16.840 0.250 17.440 ;
        RECT 24.165 16.840 25.250 17.440 ;
        RECT 39.060 16.840 40.145 17.440 ;
        RECT -0.790 16.830 0.200 16.840 ;
        RECT 24.210 16.830 25.200 16.840 ;
        RECT 39.105 16.830 40.095 16.840 ;
    END
  END vdd
  PIN vss
    ANTENNADIFFAREA 218.746887 ;
    PORT
      LAYER Pwell ;
        RECT -6.810 66.330 -5.810 69.870 ;
        RECT 60.250 68.530 60.970 69.870 ;
        RECT 60.250 66.330 61.250 68.530 ;
        RECT -6.810 58.490 -5.810 62.030 ;
        RECT 60.250 58.490 61.250 62.030 ;
        RECT -6.810 50.650 -5.810 54.190 ;
        RECT 60.250 50.650 61.250 54.190 ;
        RECT -6.810 42.810 -5.810 46.350 ;
        RECT 60.250 42.810 61.250 46.350 ;
        RECT -6.810 34.970 -5.810 38.510 ;
        RECT 60.250 34.970 61.250 38.510 ;
        RECT -6.810 27.130 -5.810 30.670 ;
        RECT 60.250 27.130 61.250 30.670 ;
        RECT -6.810 19.290 -5.810 22.830 ;
        RECT 60.250 19.290 61.250 22.830 ;
      LAYER Metal1 ;
        RECT -6.005 68.400 -5.810 69.480 ;
        RECT -6.380 67.800 -4.885 68.400 ;
        RECT 60.250 67.800 60.820 68.400 ;
        RECT -5.975 66.720 -5.810 67.800 ;
        RECT 60.250 66.720 60.445 67.800 ;
        RECT -6.005 60.560 -5.810 61.640 ;
        RECT -6.380 59.960 -5.810 60.560 ;
        RECT -6.005 58.880 -5.810 59.960 ;
        RECT 60.250 60.560 60.415 61.640 ;
        RECT 60.250 59.960 60.820 60.560 ;
        RECT 60.250 58.880 60.415 59.960 ;
        RECT -5.975 52.720 -5.810 53.800 ;
        RECT -6.380 52.120 -5.810 52.720 ;
        RECT -5.975 51.040 -5.810 52.120 ;
        RECT 60.250 52.720 60.445 53.800 ;
        RECT 60.250 52.120 60.820 52.720 ;
        RECT 60.250 51.040 60.445 52.120 ;
        RECT -6.005 44.880 -5.810 45.960 ;
        RECT -6.380 44.280 -5.810 44.880 ;
        RECT -6.005 43.200 -5.810 44.280 ;
        RECT 60.250 44.880 60.415 45.960 ;
        RECT 60.250 44.280 60.820 44.880 ;
        RECT 60.250 43.200 60.415 44.280 ;
        RECT -5.975 37.040 -5.810 38.120 ;
        RECT -6.380 36.440 -5.810 37.040 ;
        RECT -5.975 35.360 -5.810 36.440 ;
        RECT 60.250 37.040 60.445 38.120 ;
        RECT 60.250 36.440 60.820 37.040 ;
        RECT 60.250 35.360 60.445 36.440 ;
        RECT -6.005 29.200 -5.810 30.280 ;
        RECT -6.380 28.600 -5.810 29.200 ;
        RECT -6.005 27.520 -5.810 28.600 ;
        RECT 60.250 29.200 60.415 30.280 ;
        RECT 60.250 28.600 60.820 29.200 ;
        RECT 60.250 27.520 60.415 28.600 ;
        RECT -5.975 21.360 -5.810 22.440 ;
        RECT -6.380 20.760 -5.810 21.360 ;
        RECT -6.005 19.680 -5.810 20.760 ;
        RECT 60.250 21.360 60.445 22.440 ;
        RECT 60.250 20.760 60.820 21.360 ;
        RECT 60.250 19.680 60.415 20.760 ;
      LAYER Metal2 ;
        RECT 14.240 16.835 15.230 17.710 ;
        RECT 29.575 16.840 30.565 17.710 ;
        RECT 56.235 16.840 57.310 17.710 ;
    END
  END vss
  PIN reset
    ANTENNAGATEAREA 2.665600 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 60.250 66.560 60.725 66.840 ;
    END
  END reset
  PIN trim[0]
    ANTENNAGATEAREA 2.665600 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT -6.235 60.400 -5.810 60.680 ;
        RECT 60.250 60.400 60.690 60.680 ;
    END
  END trim[0]
  PIN trim[1]
    ANTENNAGATEAREA 2.665600 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT -6.250 52.560 -5.810 52.840 ;
        RECT 60.250 52.560 60.675 52.840 ;
    END
  END trim[1]
  PIN trim[2]
    ANTENNAGATEAREA 2.665600 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT -6.235 44.720 -5.810 45.000 ;
        RECT 60.250 44.720 60.690 45.000 ;
    END
  END trim[2]
  PIN trim[3]
    ANTENNAGATEAREA 2.665600 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT -6.250 36.880 -5.810 37.160 ;
        RECT 60.250 36.880 60.675 37.160 ;
    END
  END trim[3]
  PIN trim[4]
    ANTENNAGATEAREA 2.665600 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT -6.235 29.040 -5.810 29.320 ;
        RECT 60.250 29.040 60.690 29.320 ;
    END
  END trim[4]
  PIN trim[7]
    ANTENNAGATEAREA 2.665600 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT -6.235 28.480 -5.810 28.760 ;
        RECT 60.250 28.480 60.690 28.760 ;
    END
  END trim[7]
  PIN trim[8]
    ANTENNAGATEAREA 2.665600 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT -6.250 36.320 -5.810 36.600 ;
        RECT 60.250 36.320 60.690 36.600 ;
    END
  END trim[8]
  PIN trim[9]
    ANTENNAGATEAREA 2.665600 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT -6.235 44.160 -5.810 44.440 ;
        RECT 60.250 44.160 60.690 44.440 ;
    END
  END trim[9]
  PIN trim[10]
    ANTENNAGATEAREA 2.665600 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT -6.250 52.000 -5.810 52.280 ;
        RECT 60.250 52.000 60.690 52.280 ;
    END
  END trim[10]
  PIN trim[11]
    ANTENNAGATEAREA 2.665600 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT -6.235 59.840 -5.810 60.120 ;
        RECT 60.250 59.840 60.690 60.120 ;
    END
  END trim[11]
  PIN trim[12]
    ANTENNAGATEAREA 2.665600 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT -6.250 67.680 -5.810 67.960 ;
        RECT 60.250 67.680 60.705 67.960 ;
    END
  END trim[12]
  PIN trim[5]
    ANTENNAGATEAREA 2.665600 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT -6.250 21.200 -5.810 21.480 ;
        RECT 60.250 21.200 60.675 21.480 ;
    END
  END trim[5]
  PIN trim[6]
    ANTENNAGATEAREA 2.665600 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT -6.235 20.640 -5.810 20.920 ;
        RECT 60.250 20.640 60.690 20.920 ;
    END
  END trim[6]
  PIN trim[25]
    ANTENNAGATEAREA 2.665600 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT -6.250 67.120 -5.810 67.400 ;
        RECT 60.250 67.120 60.715 67.400 ;
    END
  END trim[25]
  PIN trim[13]
    ANTENNAGATEAREA 2.665600 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT -6.235 60.960 -5.810 61.240 ;
        RECT 60.250 60.960 60.690 61.240 ;
    END
  END trim[13]
  PIN trim[14]
    ANTENNAGATEAREA 2.665600 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT -6.250 53.120 -5.810 53.400 ;
        RECT 60.250 53.120 60.675 53.400 ;
    END
  END trim[14]
  PIN trim[15]
    ANTENNAGATEAREA 2.665600 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT -6.235 45.280 -5.810 45.560 ;
        RECT 60.250 45.280 60.690 45.560 ;
    END
  END trim[15]
  PIN trim[16]
    ANTENNAGATEAREA 2.665600 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT -6.250 37.440 -5.810 37.720 ;
        RECT 60.250 37.440 60.675 37.720 ;
    END
  END trim[16]
  PIN trim[17]
    ANTENNAGATEAREA 2.665600 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT -6.235 29.600 -5.810 29.880 ;
        RECT 60.250 29.600 60.690 29.880 ;
    END
  END trim[17]
  PIN trim[18]
    ANTENNAGATEAREA 2.665600 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT -6.250 21.760 -5.810 22.040 ;
        RECT 60.250 21.760 60.675 22.040 ;
    END
  END trim[18]
  PIN trim[19]
    ANTENNAGATEAREA 2.665600 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT -6.235 20.080 -5.810 20.360 ;
        RECT 60.250 20.080 60.690 20.360 ;
    END
  END trim[19]
  PIN trim[20]
    ANTENNAGATEAREA 2.665600 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT -6.235 27.920 -5.810 28.200 ;
        RECT 60.250 27.920 60.690 28.200 ;
    END
  END trim[20]
  PIN trim[21]
    ANTENNAGATEAREA 2.665600 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT -6.250 35.760 -5.810 36.040 ;
        RECT 60.250 35.760 60.675 36.040 ;
    END
  END trim[21]
  PIN trim[22]
    ANTENNAGATEAREA 2.665600 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT -6.235 43.600 -5.810 43.880 ;
        RECT 60.250 43.600 60.690 43.880 ;
    END
  END trim[22]
  PIN trim[23]
    ANTENNAGATEAREA 2.665600 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT -6.250 51.440 -5.810 51.720 ;
        RECT 60.250 51.440 60.675 51.720 ;
    END
  END trim[23]
  PIN trim[24]
    ANTENNAGATEAREA 2.665600 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT -6.235 59.280 -5.810 59.560 ;
        RECT 60.250 59.280 60.690 59.560 ;
    END
  END trim[24]
  PIN clockp[1]
    ANTENNADIFFAREA 3.712800 ;
    PORT
      LAYER Metal2 ;
        RECT 51.545 71.745 51.825 72.705 ;
    END
  END clockp[1]
  PIN clockp[0]
    ANTENNADIFFAREA 3.712800 ;
    PORT
      LAYER Metal2 ;
        RECT 43.700 71.745 43.980 72.745 ;
    END
  END clockp[0]
  OBS
      LAYER Nwell ;
        RECT -5.810 17.710 60.250 71.745 ;
      LAYER Metal1 ;
        RECT -5.810 17.710 60.250 71.745 ;
        RECT -2.370 17.670 -2.140 17.710 ;
        RECT -0.130 17.670 0.100 17.710 ;
        RECT 0.625 17.670 0.855 17.710 ;
        RECT 1.935 17.680 3.615 17.710 ;
        RECT 5.280 17.670 7.070 17.710 ;
        RECT 8.865 17.670 9.095 17.710 ;
        RECT 9.585 17.670 9.815 17.710 ;
        RECT 10.895 17.680 12.575 17.710 ;
        RECT 14.240 17.670 16.030 17.710 ;
        RECT 17.825 17.670 18.055 17.710 ;
        RECT 19.265 17.675 19.495 17.710 ;
        RECT 20.785 17.670 21.015 17.710 ;
        RECT 22.095 17.680 23.775 17.710 ;
        RECT 25.440 17.670 27.230 17.710 ;
        RECT 29.025 17.670 29.255 17.710 ;
        RECT 30.865 17.670 31.095 17.710 ;
        RECT 32.175 17.680 33.855 17.710 ;
        RECT 35.520 17.670 37.310 17.710 ;
        RECT 39.105 17.670 39.335 17.710 ;
        RECT 40.780 17.670 41.175 17.710 ;
        RECT 42.380 17.670 42.775 17.710 ;
        RECT 44.145 17.680 44.375 17.710 ;
        RECT 45.820 17.670 46.215 17.710 ;
        RECT 47.420 17.670 47.815 17.710 ;
        RECT 49.185 17.680 49.415 17.710 ;
        RECT 50.625 17.675 50.855 17.710 ;
        RECT 52.865 17.675 53.095 17.710 ;
        RECT 55.870 17.670 56.100 17.710 ;
        RECT 58.110 17.670 58.340 17.710 ;
      LAYER Metal2 ;
        RECT -4.925 17.710 59.365 71.745 ;
        RECT 28.155 17.560 28.435 17.710 ;
        RECT 32.700 17.585 32.980 17.710 ;
        RECT 40.820 17.580 41.100 17.710 ;
        RECT 50.540 17.560 50.820 17.710 ;
        RECT 28.065 17.280 28.510 17.560 ;
        RECT 50.450 17.280 50.900 17.560 ;
      LAYER Metal3 ;
        RECT -5.810 17.710 60.250 67.960 ;
        RECT 28.065 17.280 50.945 17.560 ;
  END
END ring_osc2x13
END LIBRARY

