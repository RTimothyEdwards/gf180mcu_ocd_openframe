magic
tech gf180mcuD
magscale 1 10
timestamp 1765308861
<< pwell >>
rect -364 -932 364 932
<< hvnmos >>
rect -100 -724 100 676
<< mvndiff >>
rect -188 657 -100 676
rect -188 -705 -175 657
rect -129 -705 -100 657
rect -188 -724 -100 -705
rect 100 657 188 676
rect 100 -705 129 657
rect 175 -705 188 657
rect 100 -724 188 -705
<< mvndiffc >>
rect -175 -705 -129 657
rect 129 -705 175 657
<< mvpsubdiff >>
rect -332 828 332 900
rect -332 775 -260 828
rect -332 -775 -319 775
rect -273 -775 -260 775
rect 260 775 332 828
rect -332 -828 -260 -775
rect 260 -775 273 775
rect 319 -775 332 775
rect 260 -828 332 -775
rect -332 -841 332 -828
rect -332 -887 -211 -841
rect 211 -887 332 -841
rect -332 -900 332 -887
<< mvpsubdiffcont >>
rect -319 -775 -273 775
rect 273 -775 319 775
rect -211 -887 211 -841
<< polysilicon >>
rect -100 755 100 768
rect -100 709 -70 755
rect 70 709 100 755
rect -100 676 100 709
rect -100 -768 100 -724
<< polycontact >>
rect -70 709 70 755
<< metal1 >>
rect -319 841 319 887
rect -319 775 -273 841
rect 273 775 319 841
rect -98 709 -70 755
rect 70 709 98 755
rect -175 657 -129 674
rect -175 -722 -129 -705
rect 129 657 175 674
rect 129 -722 175 -705
rect -319 -841 -273 -775
rect 273 -841 319 -775
rect -319 -887 -211 -841
rect 211 -887 319 -841
<< properties >>
string FIXED_BBOX -296 -864 296 864
string GDS_END 45276
string GDS_FILE ../gds/simple_por.gds.gz
string GDS_START 38936
<< end >>
