magic
tech gf180mcuD
magscale 1 10
timestamp 1764438222
<< metal1 >>
rect 0 133 15269 185
rect 15435 133 15452 185
rect 182 127 258 133
rect 182 101 258 110
rect 182 49 193 101
rect 245 49 258 101
rect 182 37 258 49
rect 703 127 779 133
rect 703 101 779 110
rect 703 49 715 101
rect 767 49 779 101
rect 703 37 779 49
rect 932 127 1008 133
rect 932 101 1008 110
rect 932 49 943 101
rect 995 49 1008 101
rect 932 37 1008 49
rect 1074 127 1150 133
rect 1074 101 1150 110
rect 1074 49 1085 101
rect 1137 49 1150 101
rect 1074 37 1150 49
rect 1576 127 1652 133
rect 1576 101 1652 110
rect 1576 49 1587 101
rect 1639 49 1652 101
rect 1576 37 1652 49
rect 1787 127 1863 133
rect 1787 101 1863 110
rect 1787 49 1799 101
rect 1851 49 1863 101
rect 1787 37 1863 49
rect 13244 127 13320 133
rect 13244 101 13320 110
rect 13244 49 13256 101
rect 13308 49 13320 101
rect 13244 37 13320 49
rect 13390 127 13466 133
rect 13390 101 13466 110
rect 13390 49 13402 101
rect 13454 49 13466 101
rect 13390 36 13466 49
rect 13536 127 13612 133
rect 13536 101 13612 110
rect 13536 49 13548 101
rect 13600 49 13612 101
rect 13536 37 13612 49
<< rmetal1 >>
rect 182 110 258 127
rect 703 110 779 127
rect 932 110 1008 127
rect 1074 110 1150 127
rect 1576 110 1652 127
rect 1787 110 1863 127
rect 13244 110 13320 127
rect 13390 110 13466 127
rect 13536 110 13612 127
<< via1 >>
rect 15269 133 15435 185
rect 193 49 245 101
rect 715 49 767 101
rect 943 49 995 101
rect 1085 49 1137 101
rect 1587 49 1639 101
rect 1799 49 1851 101
rect 13256 49 13308 101
rect 13402 49 13454 101
rect 13548 49 13600 101
<< metal2 >>
rect 182 101 258 232
rect 182 49 193 101
rect 245 49 258 101
rect 182 0 258 49
rect 703 101 779 232
rect 703 49 715 101
rect 767 49 779 101
rect 703 0 779 49
rect 932 101 1008 232
rect 932 49 943 101
rect 995 49 1008 101
rect 932 0 1008 49
rect 1074 101 1150 232
rect 1074 49 1085 101
rect 1137 49 1150 101
rect 1074 0 1150 49
rect 1576 101 1652 232
rect 1576 49 1587 101
rect 1639 49 1652 101
rect 1576 0 1652 49
rect 1787 101 1863 232
rect 1787 49 1799 101
rect 1851 49 1863 101
rect 1787 0 1863 49
rect 13244 101 13320 232
rect 13244 49 13256 101
rect 13308 49 13320 101
rect 13244 0 13320 49
rect 13390 101 13466 232
rect 13390 49 13402 101
rect 13454 49 13466 101
rect 13390 0 13466 49
rect 13536 101 13612 232
rect 13536 49 13548 101
rect 13600 49 13612 101
rect 13536 0 13612 49
rect 15089 0 15145 232
rect 15201 187 15257 232
rect 15201 185 15448 187
rect 15201 133 15269 185
rect 15435 133 15448 185
rect 15201 131 15448 133
rect 15201 0 15257 131
<< end >>
