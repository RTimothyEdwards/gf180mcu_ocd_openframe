magic
tech gf180mcuD
magscale 1 10
timestamp 1764438222
<< metal3 >>
rect 0 15260 303 15270
rect 0 15204 47 15260
rect 103 15204 303 15260
rect 0 15194 303 15204
rect 0 14739 303 14749
rect 0 14683 47 14739
rect 103 14683 303 14739
rect 0 14673 303 14683
rect 0 14510 303 14520
rect 0 14454 47 14510
rect 103 14454 303 14510
rect 0 14444 303 14454
rect 0 14368 303 14378
rect 0 14312 47 14368
rect 103 14312 303 14368
rect 0 14302 303 14312
rect 0 13866 303 13876
rect 0 13810 47 13866
rect 103 13810 303 13866
rect 0 13800 303 13810
rect 0 13655 303 13665
rect 0 13599 47 13655
rect 103 13599 303 13655
rect 0 13589 303 13599
rect 0 2198 303 2208
rect 0 2142 47 2198
rect 103 2142 303 2198
rect 0 2132 303 2142
rect 0 2052 303 2062
rect 0 1996 47 2052
rect 103 1996 303 2052
rect 0 1986 303 1996
rect 0 1906 303 1916
rect 0 1850 47 1906
rect 103 1850 303 1906
rect 0 1840 303 1850
rect 0 307 303 383
rect 0 182 303 251
rect 0 175 133 182
rect 189 175 303 182
rect 133 4 189 16
<< via3 >>
rect 47 15204 103 15260
rect 47 14683 103 14739
rect 47 14454 103 14510
rect 47 14312 103 14368
rect 47 13810 103 13866
rect 47 13599 103 13655
rect 47 2142 103 2198
rect 47 1996 103 2052
rect 47 1850 103 1906
rect 133 16 189 182
<< metal4 >>
rect 133 15270 189 15452
rect 37 15260 109 15270
rect 37 15204 47 15260
rect 103 15204 109 15260
rect 37 15194 109 15204
rect 125 15194 189 15270
rect 133 14749 189 15194
rect 37 14739 109 14749
rect 37 14683 47 14739
rect 103 14683 109 14739
rect 37 14673 109 14683
rect 125 14673 189 14749
rect 133 14520 189 14673
rect 37 14510 109 14520
rect 37 14454 47 14510
rect 103 14454 109 14510
rect 37 14444 109 14454
rect 125 14444 189 14520
rect 133 14378 189 14444
rect 37 14368 109 14378
rect 37 14312 47 14368
rect 103 14312 109 14368
rect 37 14302 109 14312
rect 125 14302 189 14378
rect 133 13876 189 14302
rect 37 13866 109 13876
rect 37 13810 47 13866
rect 103 13810 109 13866
rect 37 13800 109 13810
rect 125 13800 189 13876
rect 133 13665 189 13800
rect 37 13655 109 13665
rect 37 13599 47 13655
rect 103 13599 109 13655
rect 37 13589 109 13599
rect 125 13589 189 13665
rect 133 2208 189 13589
rect 37 2198 109 2208
rect 37 2142 47 2198
rect 103 2142 109 2198
rect 37 2132 109 2142
rect 125 2132 189 2208
rect 133 2062 189 2132
rect 37 2052 109 2062
rect 37 1996 47 2052
rect 103 1996 109 2052
rect 37 1986 109 1996
rect 125 1986 189 2062
rect 133 1916 189 1986
rect 37 1906 109 1916
rect 37 1850 47 1906
rect 103 1850 109 1906
rect 37 1840 109 1850
rect 125 1840 189 1916
rect 133 182 189 1840
rect 133 0 189 16
<< rmetal4 >>
rect 109 15194 125 15270
rect 109 14673 125 14749
rect 109 14444 125 14520
rect 109 14302 125 14378
rect 109 13800 125 13876
rect 109 13589 125 13665
rect 109 2132 125 2208
rect 109 1986 125 2062
rect 109 1840 125 1916
<< properties >>
string flatten true
<< end >>
