magic
tech gf180mcuD
magscale 1 10
timestamp 1764176821
<< metal2 >>
rect 0 14444 271 14456
rect 0 12568 2 14444
rect 269 12568 271 14444
rect 0 12556 271 12568
rect 0 11964 271 11976
rect 0 9938 2 11964
rect 269 9938 271 11964
rect 0 9926 271 9938
rect 0 9594 271 9606
rect 0 7568 2 9594
rect 269 7568 271 9594
rect 0 7556 271 7568
rect 0 6888 271 6900
rect 0 4862 2 6888
rect 269 4862 271 6888
rect 0 4850 271 4862
rect 0 4518 271 4530
rect 0 2492 2 4518
rect 269 2492 271 4518
rect 0 2480 271 2492
rect 0 1888 271 1900
rect 0 12 2 1888
rect 269 12 271 1888
rect 0 0 271 12
<< via2 >>
rect 2 12568 269 14444
rect 2 9938 269 11964
rect 2 7568 269 9594
rect 2 4862 269 6888
rect 2 2492 269 4518
rect 2 12 269 1888
<< metal3 >>
rect 0 14444 271 14456
rect 0 12568 2 14444
rect 269 12568 271 14444
rect 0 11964 271 12568
rect 0 9938 2 11964
rect 269 9938 271 11964
rect 0 9594 271 9938
rect 0 7568 2 9594
rect 269 7568 271 9594
rect 0 6888 271 7568
rect 0 4862 2 6888
rect 269 4862 271 6888
rect 0 4518 271 4862
rect 0 2492 2 4518
rect 269 2492 271 4518
rect 0 1888 271 2492
rect 0 12 2 1888
rect 269 12 271 1888
rect 0 0 271 12
<< via3 >>
rect 2 12568 269 14444
rect 2 9938 269 11964
rect 2 7568 269 9594
rect 2 4862 269 6888
rect 2 2492 269 4518
rect 2 12 269 1888
<< metal4 >>
rect 0 14444 271 14456
rect 0 12568 2 14444
rect 269 12568 271 14444
rect 0 12556 271 12568
rect 0 11964 271 11976
rect 0 9938 2 11964
rect 269 9938 271 11964
rect 0 9926 271 9938
rect 0 9594 271 9606
rect 0 7568 2 9594
rect 269 7568 271 9594
rect 0 7556 271 7568
rect 0 6888 271 6900
rect 0 4862 2 6888
rect 269 4862 271 6888
rect 0 4850 271 4862
rect 0 4518 271 4530
rect 0 2492 2 4518
rect 269 2492 271 4518
rect 0 2480 271 2492
rect 0 1888 271 1900
rect 0 12 2 1888
rect 269 12 271 1888
rect 0 0 271 12
<< via4 >>
rect 2 12568 269 14444
rect 2 9938 269 11964
rect 2 7568 269 9594
rect 2 4862 269 6888
rect 2 2492 269 4518
rect 2 12 269 1888
<< metal5 >>
rect 0 14444 271 14456
rect 0 12568 2 14444
rect 269 12568 271 14444
rect 0 12556 271 12568
rect 0 11964 271 11976
rect 0 9938 2 11964
rect 269 9938 271 11964
rect 0 9926 271 9938
rect 0 9594 271 9606
rect 0 7568 2 9594
rect 269 7568 271 9594
rect 0 7556 271 7568
rect 0 6888 271 6900
rect 0 4862 2 6888
rect 269 4862 271 6888
rect 0 4850 271 4862
rect 0 4518 271 4530
rect 0 2492 2 4518
rect 269 2492 271 4518
rect 0 2480 271 2492
rect 0 1888 271 1900
rect 0 12 2 1888
rect 269 12 271 1888
rect 0 0 271 12
<< properties >>
string flatten true
<< end >>
