magic
tech gf180mcuD
magscale 1 10
timestamp 1765305544
<< error_p >>
rect 528544 136422 528554 136432
rect 528932 136422 528942 136432
rect 539544 136426 539554 136436
rect 539934 136426 539944 136436
rect 550544 136426 550554 136436
rect 550934 136426 550944 136436
rect 561544 136426 561554 136436
rect 561934 136426 561944 136436
rect 572544 136426 572554 136436
rect 572934 136426 572944 136436
rect 528534 136412 528544 136422
rect 528942 136412 528952 136422
rect 539534 136416 539544 136426
rect 539944 136416 539954 136426
rect 550534 136416 550544 136426
rect 550944 136416 550954 136426
rect 561534 136416 561544 136426
rect 561944 136416 561954 136426
rect 572534 136416 572544 136426
rect 572944 136416 572954 136426
rect 583544 136422 583554 136432
rect 583934 136422 583944 136432
rect 583534 136412 583544 136422
rect 583944 136412 583954 136422
rect 528534 135728 528544 135738
rect 528942 135728 528952 135738
rect 539534 135729 539544 135739
rect 539944 135729 539954 135739
rect 528544 135718 528554 135728
rect 528932 135718 528942 135728
rect 539544 135719 539554 135729
rect 539934 135719 539944 135729
rect 550534 135726 550544 135736
rect 550944 135726 550954 135736
rect 561534 135726 561544 135736
rect 561944 135726 561954 135736
rect 572534 135727 572544 135737
rect 572944 135727 572954 135737
rect 550544 135716 550554 135726
rect 550934 135716 550944 135726
rect 561544 135716 561554 135726
rect 561934 135716 561944 135726
rect 572544 135717 572554 135727
rect 572934 135717 572944 135727
rect 583534 135726 583544 135736
rect 583944 135726 583954 135736
rect 583544 135716 583554 135726
rect 583934 135716 583944 135726
rect 573284 135547 573294 135557
rect 573674 135547 573684 135557
rect 584284 135547 584294 135557
rect 584674 135547 584684 135557
rect 573274 135537 573284 135547
rect 573684 135537 573694 135547
rect 584274 135537 584284 135547
rect 584684 135537 584694 135547
rect 529284 135510 529294 135520
rect 529674 135510 529684 135520
rect 540284 135510 540294 135520
rect 540674 135510 540684 135520
rect 529274 135500 529284 135510
rect 529684 135500 529694 135510
rect 540274 135500 540284 135510
rect 540684 135500 540694 135510
rect 573274 135337 573284 135347
rect 573684 135337 573694 135347
rect 584274 135337 584284 135347
rect 584684 135337 584694 135347
rect 573284 135327 573294 135337
rect 573674 135327 573684 135337
rect 584284 135327 584294 135337
rect 584674 135327 584684 135337
rect 529274 135300 529284 135310
rect 529684 135300 529694 135310
rect 540274 135300 540284 135310
rect 540684 135300 540694 135310
rect 529284 135290 529294 135300
rect 529674 135290 529684 135300
rect 540284 135290 540294 135300
rect 540674 135290 540684 135300
rect 573284 134335 573294 134345
rect 573674 134335 573684 134345
rect 584284 134335 584294 134345
rect 584674 134335 584684 134345
rect 573274 134325 573284 134335
rect 573684 134325 573694 134335
rect 584274 134325 584284 134335
rect 584684 134325 584694 134335
rect 529284 134298 529294 134308
rect 529674 134298 529684 134308
rect 540284 134298 540294 134308
rect 540674 134298 540684 134308
rect 529274 134288 529284 134298
rect 529684 134288 529694 134298
rect 540274 134288 540284 134298
rect 540684 134288 540694 134298
rect 573274 134125 573284 134135
rect 573684 134125 573694 134135
rect 584274 134125 584284 134135
rect 584684 134125 584694 134135
rect 573284 134115 573294 134125
rect 573674 134115 573684 134125
rect 584284 134115 584294 134125
rect 584674 134115 584684 134125
rect 529274 134088 529284 134098
rect 529684 134088 529694 134098
rect 540274 134088 540284 134098
rect 540684 134088 540694 134098
rect 529284 134078 529294 134088
rect 529674 134078 529684 134088
rect 540284 134078 540294 134088
rect 540674 134078 540684 134088
rect 573284 133123 573294 133133
rect 573674 133123 573684 133133
rect 584284 133123 584294 133133
rect 584674 133123 584684 133133
rect 573274 133113 573284 133123
rect 573684 133113 573694 133123
rect 584274 133113 584284 133123
rect 584684 133113 584694 133123
rect 529284 133086 529294 133096
rect 529674 133086 529684 133096
rect 540284 133086 540294 133096
rect 540674 133086 540684 133096
rect 529274 133076 529284 133086
rect 529684 133076 529694 133086
rect 540274 133076 540284 133086
rect 540684 133076 540694 133086
rect 573274 132913 573284 132923
rect 573684 132913 573694 132923
rect 584274 132913 584284 132923
rect 584684 132913 584694 132923
rect 573284 132903 573294 132913
rect 573674 132903 573684 132913
rect 584284 132903 584294 132913
rect 584674 132903 584684 132913
rect 529274 132876 529284 132886
rect 529684 132876 529694 132886
rect 540274 132876 540284 132886
rect 540684 132876 540694 132886
rect 529284 132866 529294 132876
rect 529674 132866 529684 132876
rect 540284 132866 540294 132876
rect 540674 132866 540684 132876
rect 573284 131911 573294 131921
rect 573674 131911 573684 131921
rect 584284 131911 584294 131921
rect 584674 131911 584684 131921
rect 573274 131901 573284 131911
rect 573684 131901 573694 131911
rect 584274 131901 584284 131911
rect 584684 131901 584694 131911
rect 529284 131874 529294 131884
rect 529674 131874 529684 131884
rect 540284 131874 540294 131884
rect 540674 131874 540684 131884
rect 529274 131864 529284 131874
rect 529684 131864 529694 131874
rect 540274 131864 540284 131874
rect 540684 131864 540694 131874
rect 573274 131701 573284 131711
rect 573684 131701 573694 131711
rect 584274 131701 584284 131711
rect 584684 131701 584694 131711
rect 573284 131691 573294 131701
rect 573674 131691 573684 131701
rect 584284 131691 584294 131701
rect 584674 131691 584684 131701
rect 529274 131664 529284 131674
rect 529684 131664 529694 131674
rect 540274 131664 540284 131674
rect 540684 131664 540694 131674
rect 529284 131654 529294 131664
rect 529674 131654 529684 131664
rect 540284 131654 540294 131664
rect 540674 131654 540684 131664
rect 573284 130699 573294 130709
rect 573674 130699 573684 130709
rect 584284 130699 584294 130709
rect 584674 130699 584684 130709
rect 573274 130689 573284 130699
rect 573684 130689 573694 130699
rect 584274 130689 584284 130699
rect 584684 130689 584694 130699
rect 529284 130662 529294 130672
rect 529674 130662 529684 130672
rect 540284 130662 540294 130672
rect 540674 130662 540684 130672
rect 529274 130652 529284 130662
rect 529684 130652 529694 130662
rect 540274 130652 540284 130662
rect 540684 130652 540694 130662
rect 573274 130489 573284 130499
rect 573684 130489 573694 130499
rect 584274 130489 584284 130499
rect 584684 130489 584694 130499
rect 573284 130479 573294 130489
rect 573674 130479 573684 130489
rect 584284 130479 584294 130489
rect 584674 130479 584684 130489
rect 529274 130452 529284 130462
rect 529684 130452 529694 130462
rect 540274 130452 540284 130462
rect 540684 130452 540694 130462
rect 529284 130442 529294 130452
rect 529674 130442 529684 130452
rect 540284 130442 540294 130452
rect 540674 130442 540684 130452
rect 573284 129487 573294 129497
rect 573674 129487 573684 129497
rect 584284 129487 584294 129497
rect 584674 129487 584684 129497
rect 573274 129477 573284 129487
rect 573684 129477 573694 129487
rect 584274 129477 584284 129487
rect 584684 129477 584694 129487
rect 529284 129450 529294 129460
rect 529674 129450 529684 129460
rect 540284 129450 540294 129460
rect 540674 129450 540684 129460
rect 529274 129440 529284 129450
rect 529684 129440 529694 129450
rect 540274 129440 540284 129450
rect 540684 129440 540694 129450
rect 573274 129277 573284 129287
rect 573684 129277 573694 129287
rect 584274 129277 584284 129287
rect 584684 129277 584694 129287
rect 573284 129267 573294 129277
rect 573674 129267 573684 129277
rect 584284 129267 584294 129277
rect 584674 129267 584684 129277
rect 529274 129240 529284 129250
rect 529684 129240 529694 129250
rect 540274 129240 540284 129250
rect 540684 129240 540694 129250
rect 529284 129230 529294 129240
rect 529674 129230 529684 129240
rect 540284 129230 540294 129240
rect 540674 129230 540684 129240
rect 573284 128275 573294 128285
rect 573674 128275 573684 128285
rect 584284 128275 584294 128285
rect 584674 128275 584684 128285
rect 573274 128265 573284 128275
rect 573684 128265 573694 128275
rect 584274 128265 584284 128275
rect 584684 128265 584694 128275
rect 529284 128238 529294 128248
rect 529674 128238 529684 128248
rect 540284 128238 540294 128248
rect 540674 128238 540684 128248
rect 529274 128228 529284 128238
rect 529684 128228 529694 128238
rect 540274 128228 540284 128238
rect 540684 128228 540694 128238
rect 573274 128065 573284 128075
rect 573684 128065 573694 128075
rect 584274 128065 584284 128075
rect 584684 128065 584694 128075
rect 573284 128055 573294 128065
rect 573674 128055 573684 128065
rect 584284 128055 584294 128065
rect 584674 128055 584684 128065
rect 529274 128028 529284 128038
rect 529684 128028 529694 128038
rect 540274 128028 540284 128038
rect 540684 128028 540694 128038
rect 529284 128018 529294 128028
rect 529674 128018 529684 128028
rect 540284 128018 540294 128028
rect 540674 128018 540684 128028
rect 573284 127063 573294 127073
rect 573674 127063 573684 127073
rect 584284 127063 584294 127073
rect 584674 127063 584684 127073
rect 573274 127053 573284 127063
rect 573684 127053 573694 127063
rect 584274 127053 584284 127063
rect 584684 127053 584694 127063
rect 529284 127026 529294 127036
rect 529674 127026 529684 127036
rect 540284 127026 540294 127036
rect 540674 127026 540684 127036
rect 529274 127016 529284 127026
rect 529684 127016 529694 127026
rect 540274 127016 540284 127026
rect 540684 127016 540694 127026
rect 573274 126853 573284 126863
rect 573684 126853 573694 126863
rect 584274 126853 584284 126863
rect 584684 126853 584694 126863
rect 573284 126843 573294 126853
rect 573674 126843 573684 126853
rect 584284 126843 584294 126853
rect 584674 126843 584684 126853
rect 529274 126816 529284 126826
rect 529684 126816 529694 126826
rect 540274 126816 540284 126826
rect 540684 126816 540694 126826
rect 529284 126806 529294 126816
rect 529674 126806 529684 126816
rect 540284 126806 540294 126816
rect 540674 126806 540684 126816
rect 573284 125851 573294 125861
rect 573674 125851 573684 125861
rect 584284 125851 584294 125861
rect 584674 125851 584684 125861
rect 573274 125841 573284 125851
rect 573684 125841 573694 125851
rect 584274 125841 584284 125851
rect 584684 125841 584694 125851
rect 529284 125814 529294 125824
rect 529674 125814 529684 125824
rect 540284 125814 540294 125824
rect 540674 125814 540684 125824
rect 529274 125804 529284 125814
rect 529684 125804 529694 125814
rect 540274 125804 540284 125814
rect 540684 125804 540694 125814
rect 573274 125641 573284 125651
rect 573684 125641 573694 125651
rect 584274 125641 584284 125651
rect 584684 125641 584694 125651
rect 573284 125631 573294 125641
rect 573674 125631 573684 125641
rect 584284 125631 584294 125641
rect 584674 125631 584684 125641
rect 529274 125604 529284 125614
rect 529684 125604 529694 125614
rect 540274 125604 540284 125614
rect 540684 125604 540694 125614
rect 529284 125594 529294 125604
rect 529674 125594 529684 125604
rect 540284 125594 540294 125604
rect 540674 125594 540684 125604
rect 573284 124639 573294 124649
rect 573674 124639 573684 124649
rect 584284 124639 584294 124649
rect 584674 124639 584684 124649
rect 573274 124629 573284 124639
rect 573684 124629 573694 124639
rect 584274 124629 584284 124639
rect 584684 124629 584694 124639
rect 529284 124602 529294 124612
rect 529674 124602 529684 124612
rect 540284 124602 540294 124612
rect 540674 124602 540684 124612
rect 529274 124592 529284 124602
rect 529684 124592 529694 124602
rect 540274 124592 540284 124602
rect 540684 124592 540694 124602
rect 573274 124429 573284 124439
rect 573684 124429 573694 124439
rect 584274 124429 584284 124439
rect 584684 124429 584694 124439
rect 573284 124419 573294 124429
rect 573674 124419 573684 124429
rect 584284 124419 584294 124429
rect 584674 124419 584684 124429
rect 529274 124392 529284 124402
rect 529684 124392 529694 124402
rect 540274 124392 540284 124402
rect 540684 124392 540694 124402
rect 529284 124382 529294 124392
rect 529674 124382 529684 124392
rect 540284 124382 540294 124392
rect 540674 124382 540684 124392
rect 573284 123427 573294 123437
rect 573674 123427 573684 123437
rect 584284 123427 584294 123437
rect 584674 123427 584684 123437
rect 573274 123417 573284 123427
rect 573684 123417 573694 123427
rect 584274 123417 584284 123427
rect 584684 123417 584694 123427
rect 529284 123390 529294 123400
rect 529674 123390 529684 123400
rect 540284 123390 540294 123400
rect 540674 123390 540684 123400
rect 529274 123380 529284 123390
rect 529684 123380 529694 123390
rect 540274 123380 540284 123390
rect 540684 123380 540694 123390
rect 573274 123217 573284 123227
rect 573684 123217 573694 123227
rect 584274 123217 584284 123227
rect 584684 123217 584694 123227
rect 573284 123207 573294 123217
rect 573674 123207 573684 123217
rect 584284 123207 584294 123217
rect 584674 123207 584684 123217
rect 529274 123180 529284 123190
rect 529684 123180 529694 123190
rect 540274 123180 540284 123190
rect 540684 123180 540694 123190
rect 529284 123170 529294 123180
rect 529674 123170 529684 123180
rect 540284 123170 540294 123180
rect 540674 123170 540684 123180
rect 573284 122215 573294 122225
rect 573674 122215 573684 122225
rect 584284 122215 584294 122225
rect 584674 122215 584684 122225
rect 573274 122205 573284 122215
rect 573684 122205 573694 122215
rect 584274 122205 584284 122215
rect 584684 122205 584694 122215
rect 529284 122178 529294 122188
rect 529674 122178 529684 122188
rect 540284 122178 540294 122188
rect 540674 122178 540684 122188
rect 529274 122168 529284 122178
rect 529684 122168 529694 122178
rect 540274 122168 540284 122178
rect 540684 122168 540694 122178
rect 573274 122005 573284 122015
rect 573684 122005 573694 122015
rect 584274 122005 584284 122015
rect 584684 122005 584694 122015
rect 573284 121995 573294 122005
rect 573674 121995 573684 122005
rect 584284 121995 584294 122005
rect 584674 121995 584684 122005
rect 529274 121968 529284 121978
rect 529684 121968 529694 121978
rect 540274 121968 540284 121978
rect 540684 121968 540694 121978
rect 529284 121958 529294 121968
rect 529674 121958 529684 121968
rect 540284 121958 540294 121968
rect 540674 121958 540684 121968
rect 573284 121003 573294 121013
rect 573674 121003 573684 121013
rect 584284 121003 584294 121013
rect 584674 121003 584684 121013
rect 573274 120993 573284 121003
rect 573684 120993 573694 121003
rect 584274 120993 584284 121003
rect 584684 120993 584694 121003
rect 529284 120966 529294 120976
rect 529674 120966 529684 120976
rect 540284 120966 540294 120976
rect 540674 120966 540684 120976
rect 529274 120956 529284 120966
rect 529684 120956 529694 120966
rect 540274 120956 540284 120966
rect 540684 120956 540694 120966
rect 573274 120793 573284 120803
rect 573684 120793 573694 120803
rect 584274 120793 584284 120803
rect 584684 120793 584694 120803
rect 573284 120783 573294 120793
rect 573674 120783 573684 120793
rect 584284 120783 584294 120793
rect 584674 120783 584684 120793
rect 529274 120756 529284 120766
rect 529684 120756 529694 120766
rect 540274 120756 540284 120766
rect 540684 120756 540694 120766
rect 529284 120746 529294 120756
rect 529674 120746 529684 120756
rect 540284 120746 540294 120756
rect 540674 120746 540684 120756
rect 573284 119791 573294 119801
rect 573674 119791 573684 119801
rect 584284 119791 584294 119801
rect 584674 119791 584684 119801
rect 573274 119781 573284 119791
rect 573684 119781 573694 119791
rect 584274 119781 584284 119791
rect 584684 119781 584694 119791
rect 529284 119754 529294 119764
rect 529674 119754 529684 119764
rect 540284 119754 540294 119764
rect 540674 119754 540684 119764
rect 529274 119744 529284 119754
rect 529684 119744 529694 119754
rect 540274 119744 540284 119754
rect 540684 119744 540694 119754
rect 573274 119581 573284 119591
rect 573684 119581 573694 119591
rect 584274 119581 584284 119591
rect 584684 119581 584694 119591
rect 573284 119571 573294 119581
rect 573674 119571 573684 119581
rect 584284 119571 584294 119581
rect 584674 119571 584684 119581
rect 529274 119544 529284 119554
rect 529684 119544 529694 119554
rect 540274 119544 540284 119554
rect 540684 119544 540694 119554
rect 529284 119534 529294 119544
rect 529674 119534 529684 119544
rect 540284 119534 540294 119544
rect 540674 119534 540684 119544
rect 573284 118579 573294 118589
rect 573674 118579 573684 118589
rect 584284 118579 584294 118589
rect 584674 118579 584684 118589
rect 573274 118569 573284 118579
rect 573684 118569 573694 118579
rect 584274 118569 584284 118579
rect 584684 118569 584694 118579
rect 529284 118542 529294 118552
rect 529674 118542 529684 118552
rect 540284 118542 540294 118552
rect 540674 118542 540684 118552
rect 529274 118532 529284 118542
rect 529684 118532 529694 118542
rect 540274 118532 540284 118542
rect 540684 118532 540694 118542
rect 573274 118369 573284 118379
rect 573684 118369 573694 118379
rect 584274 118369 584284 118379
rect 584684 118369 584694 118379
rect 573284 118359 573294 118369
rect 573674 118359 573684 118369
rect 584284 118359 584294 118369
rect 584674 118359 584684 118369
rect 529274 118332 529284 118342
rect 529684 118332 529694 118342
rect 540274 118332 540284 118342
rect 540684 118332 540694 118342
rect 529284 118322 529294 118332
rect 529674 118322 529684 118332
rect 540284 118322 540294 118332
rect 540674 118322 540684 118332
rect 573284 117367 573294 117377
rect 573674 117367 573684 117377
rect 584284 117367 584294 117377
rect 584674 117367 584684 117377
rect 573274 117357 573284 117367
rect 573684 117357 573694 117367
rect 584274 117357 584284 117367
rect 584684 117357 584694 117367
rect 529284 117330 529294 117340
rect 529674 117330 529684 117340
rect 540284 117330 540294 117340
rect 540674 117330 540684 117340
rect 529274 117320 529284 117330
rect 529684 117320 529694 117330
rect 540274 117320 540284 117330
rect 540684 117320 540694 117330
rect 573274 117157 573284 117167
rect 573684 117157 573694 117167
rect 584274 117157 584284 117167
rect 584684 117157 584694 117167
rect 573284 117147 573294 117157
rect 573674 117147 573684 117157
rect 584284 117147 584294 117157
rect 584674 117147 584684 117157
rect 529274 117120 529284 117130
rect 529684 117120 529694 117130
rect 540274 117120 540284 117130
rect 540684 117120 540694 117130
rect 529284 117110 529294 117120
rect 529674 117110 529684 117120
rect 540284 117110 540294 117120
rect 540674 117110 540684 117120
rect 573284 116155 573294 116165
rect 573674 116155 573684 116165
rect 584284 116155 584294 116165
rect 584674 116155 584684 116165
rect 573274 116145 573284 116155
rect 573684 116145 573694 116155
rect 584274 116145 584284 116155
rect 584684 116145 584694 116155
rect 529284 116118 529294 116128
rect 529674 116118 529684 116128
rect 540284 116118 540294 116128
rect 540674 116118 540684 116128
rect 529274 116108 529284 116118
rect 529684 116108 529694 116118
rect 540274 116108 540284 116118
rect 540684 116108 540694 116118
rect 573274 115945 573284 115955
rect 573684 115945 573694 115955
rect 584274 115945 584284 115955
rect 584684 115945 584694 115955
rect 573284 115935 573294 115945
rect 573674 115935 573684 115945
rect 584284 115935 584294 115945
rect 584674 115935 584684 115945
rect 529274 115908 529284 115918
rect 529684 115908 529694 115918
rect 540274 115908 540284 115918
rect 540684 115908 540694 115918
rect 529284 115898 529294 115908
rect 529674 115898 529684 115908
rect 540284 115898 540294 115908
rect 540674 115898 540684 115908
rect 529284 114875 529294 114885
rect 529674 114875 529684 114885
rect 540284 114875 540294 114885
rect 540674 114875 540684 114885
rect 573284 114880 573294 114890
rect 573674 114880 573684 114890
rect 529274 114865 529284 114875
rect 529684 114865 529694 114875
rect 540274 114865 540284 114875
rect 540684 114865 540694 114875
rect 573274 114870 573284 114880
rect 573684 114870 573694 114880
rect 584284 114875 584294 114885
rect 584674 114875 584684 114885
rect 584274 114865 584284 114875
rect 584684 114865 584694 114875
rect 573274 114727 573284 114737
rect 573684 114727 573694 114737
rect 573284 114717 573294 114727
rect 573674 114717 573684 114727
rect 584274 114725 584284 114735
rect 584684 114725 584694 114735
rect 584284 114715 584294 114725
rect 584674 114715 584684 114725
rect 529274 114675 529284 114685
rect 529684 114675 529694 114685
rect 540274 114675 540284 114685
rect 540684 114675 540694 114685
rect 529284 114665 529294 114675
rect 529674 114665 529684 114675
rect 540284 114665 540294 114675
rect 540674 114665 540684 114675
rect 529284 114606 529294 114616
rect 529674 114606 529684 114616
rect 540284 114606 540294 114616
rect 540674 114606 540684 114616
rect 529274 114596 529284 114606
rect 529684 114596 529694 114606
rect 540274 114596 540284 114606
rect 540684 114596 540694 114606
rect 573284 114604 573294 114614
rect 573674 114604 573684 114614
rect 584284 114605 584294 114615
rect 584674 114605 584684 114615
rect 573274 114594 573284 114604
rect 573684 114594 573694 114604
rect 584274 114595 584284 114605
rect 584684 114595 584694 114605
rect 529274 114270 529284 114280
rect 529684 114270 529694 114280
rect 540274 114270 540284 114280
rect 540684 114270 540694 114280
rect 573274 114270 573284 114280
rect 573684 114270 573694 114280
rect 584274 114270 584284 114280
rect 584684 114270 584694 114280
rect 529284 114260 529294 114270
rect 529674 114260 529684 114270
rect 540284 114260 540294 114270
rect 540674 114260 540684 114270
rect 573284 114260 573294 114270
rect 573674 114260 573684 114270
rect 584284 114260 584294 114270
rect 584674 114260 584684 114270
rect 528544 113982 528554 113992
rect 528934 113982 528944 113992
rect 539544 113982 539554 113992
rect 539934 113982 539944 113992
rect 528534 113972 528544 113982
rect 528944 113972 528954 113982
rect 539534 113972 539544 113982
rect 539944 113972 539954 113982
rect 572544 113978 572554 113988
rect 572934 113978 572944 113988
rect 583544 113981 583554 113991
rect 583934 113981 583944 113991
rect 572534 113968 572544 113978
rect 572944 113968 572954 113978
rect 583534 113971 583544 113981
rect 583944 113971 583954 113981
rect 550544 112764 550554 112774
rect 550934 112764 550944 112774
rect 561544 112764 561554 112774
rect 561934 112764 561944 112774
rect 550534 112754 550544 112764
rect 550944 112754 550954 112764
rect 561534 112754 561544 112764
rect 561944 112754 561954 112764
rect 528534 112576 528544 112586
rect 528944 112576 528954 112586
rect 539534 112576 539544 112586
rect 539944 112576 539954 112586
rect 572534 112585 572544 112595
rect 572944 112585 572954 112595
rect 528544 112566 528554 112576
rect 528934 112566 528944 112576
rect 539544 112566 539554 112576
rect 539934 112566 539944 112576
rect 572544 112575 572554 112585
rect 572934 112575 572944 112585
rect 583534 112577 583544 112587
rect 583944 112577 583954 112587
rect 583544 112567 583554 112577
rect 583934 112567 583944 112577
rect 550534 112303 550544 112313
rect 550944 112303 550954 112313
rect 561534 112303 561544 112313
rect 561944 112303 561954 112313
rect 550544 112293 550554 112303
rect 550934 112293 550944 112303
rect 561544 112293 561554 112303
rect 561934 112293 561944 112303
rect 550544 111567 550554 111577
rect 550934 111567 550944 111577
rect 550534 111557 550544 111567
rect 550944 111557 550954 111567
rect 561544 111562 561554 111572
rect 561934 111562 561944 111572
rect 561534 111552 561544 111562
rect 561944 111552 561954 111562
rect 528544 111234 528554 111244
rect 528934 111234 528944 111244
rect 583544 111234 583554 111244
rect 583934 111234 583944 111244
rect 528534 111224 528544 111234
rect 528944 111224 528954 111234
rect 583534 111224 583544 111234
rect 583944 111224 583954 111234
rect 528534 111035 528544 111045
rect 528944 111035 528954 111045
rect 583534 111036 583544 111046
rect 583944 111036 583954 111046
rect 528544 111025 528554 111035
rect 528934 111025 528944 111035
rect 583544 111026 583554 111036
rect 583934 111026 583944 111036
rect 529284 110765 529294 110775
rect 529674 110765 529684 110775
rect 540284 110765 540294 110775
rect 540674 110765 540684 110775
rect 573284 110765 573294 110775
rect 573674 110765 573684 110775
rect 584284 110765 584294 110775
rect 584674 110765 584684 110775
rect 529274 110755 529284 110765
rect 529684 110755 529694 110765
rect 540274 110755 540284 110765
rect 540684 110755 540694 110765
rect 573274 110755 573284 110765
rect 573684 110755 573694 110765
rect 584274 110755 584284 110765
rect 584684 110755 584694 110765
rect 550534 110083 550544 110093
rect 550944 110083 550954 110093
rect 561534 110084 561544 110094
rect 561944 110084 561954 110094
rect 550544 110073 550554 110083
rect 550934 110073 550944 110083
rect 561544 110074 561554 110084
rect 561934 110074 561944 110084
rect 529274 109365 529284 109375
rect 529684 109365 529694 109375
rect 540274 109365 540284 109375
rect 540684 109365 540694 109375
rect 573274 109365 573284 109375
rect 573684 109365 573694 109375
rect 584274 109366 584284 109376
rect 584684 109366 584694 109376
rect 529284 109355 529294 109365
rect 529674 109355 529684 109365
rect 540284 109355 540294 109365
rect 540674 109355 540684 109365
rect 573284 109355 573294 109365
rect 573674 109355 573684 109365
rect 584284 109356 584294 109366
rect 584674 109356 584684 109366
rect 539544 107290 539554 107300
rect 539934 107290 539944 107300
rect 572544 107290 572554 107300
rect 572934 107290 572944 107300
rect 583544 107290 583554 107300
rect 583934 107290 583944 107300
rect 528544 107280 528554 107290
rect 528934 107280 528944 107290
rect 539534 107280 539544 107290
rect 539944 107280 539954 107290
rect 572534 107280 572544 107290
rect 572944 107280 572954 107290
rect 583534 107280 583544 107290
rect 583944 107280 583954 107290
rect 528534 107270 528544 107280
rect 528944 107270 528954 107280
rect 528534 106971 528544 106981
rect 528944 106971 528954 106981
rect 528544 106961 528554 106971
rect 528934 106961 528944 106971
rect 583534 106906 583544 106916
rect 583944 106906 583954 106916
rect 583544 106896 583554 106906
rect 583934 106896 583944 106906
rect 539534 106848 539544 106858
rect 539944 106848 539954 106858
rect 572534 106848 572544 106858
rect 572944 106848 572954 106858
rect 539544 106838 539554 106848
rect 539934 106838 539944 106848
rect 572544 106838 572554 106848
rect 572934 106838 572944 106848
rect 529284 106702 529294 106712
rect 529674 106702 529684 106712
rect 540284 106702 540294 106712
rect 540674 106702 540684 106712
rect 573284 106702 573294 106712
rect 573674 106702 573684 106712
rect 584284 106702 584294 106712
rect 584674 106702 584684 106712
rect 529274 106692 529284 106702
rect 529684 106692 529694 106702
rect 540274 106692 540284 106702
rect 540684 106692 540694 106702
rect 573274 106692 573284 106702
rect 573684 106692 573694 106702
rect 584274 106692 584284 106702
rect 584684 106692 584694 106702
rect 540274 106270 540284 106280
rect 540684 106270 540694 106280
rect 573274 106270 573284 106280
rect 573684 106270 573694 106280
rect 529274 106253 529284 106263
rect 529684 106253 529694 106263
rect 540284 106260 540294 106270
rect 540674 106260 540684 106270
rect 573284 106260 573294 106270
rect 573674 106260 573684 106270
rect 584274 106256 584284 106266
rect 584684 106256 584694 106266
rect 529284 106243 529294 106253
rect 529674 106243 529684 106253
rect 584284 106246 584294 106256
rect 584674 106246 584684 106256
rect 528544 105548 528554 105558
rect 528934 105548 528944 105558
rect 539544 105552 539554 105562
rect 539934 105552 539944 105562
rect 572544 105552 572554 105562
rect 572934 105552 572944 105562
rect 583544 105552 583554 105562
rect 583934 105552 583944 105562
rect 528534 105538 528544 105548
rect 528944 105538 528954 105548
rect 539534 105542 539544 105552
rect 539944 105542 539954 105552
rect 572534 105542 572544 105552
rect 572944 105542 572954 105552
rect 583534 105542 583544 105552
rect 583944 105542 583954 105552
rect 528534 103642 528544 103652
rect 528944 103642 528954 103652
rect 539534 103645 539544 103655
rect 539944 103645 539954 103655
rect 572534 103645 572544 103655
rect 572944 103645 572954 103655
rect 583534 103645 583544 103655
rect 583944 103645 583954 103655
rect 528544 103632 528554 103642
rect 528934 103632 528944 103642
rect 539544 103635 539554 103645
rect 539934 103635 539944 103645
rect 572544 103635 572554 103645
rect 572934 103635 572944 103645
rect 583544 103635 583554 103645
rect 583934 103635 583944 103645
rect 529284 103445 529294 103455
rect 529674 103445 529684 103455
rect 540284 103445 540294 103455
rect 540674 103445 540684 103455
rect 529274 103435 529284 103445
rect 529684 103435 529694 103445
rect 540274 103435 540284 103445
rect 540684 103435 540694 103445
rect 573284 103441 573294 103451
rect 573674 103441 573684 103451
rect 584284 103445 584294 103455
rect 584674 103445 584684 103455
rect 573274 103431 573284 103441
rect 573684 103431 573694 103441
rect 584274 103435 584284 103445
rect 584684 103435 584694 103445
rect 529274 101588 529284 101598
rect 529684 101588 529694 101598
rect 540274 101588 540284 101598
rect 540684 101588 540694 101598
rect 573274 101588 573284 101598
rect 573684 101588 573694 101598
rect 584274 101589 584284 101599
rect 584684 101589 584694 101599
rect 529284 101578 529294 101588
rect 529674 101578 529684 101588
rect 540284 101578 540294 101588
rect 540674 101578 540684 101588
rect 573284 101578 573294 101588
rect 573674 101578 573684 101588
rect 584284 101579 584294 101589
rect 584674 101579 584684 101589
rect 528544 101463 528554 101473
rect 528934 101463 528944 101473
rect 528534 101453 528544 101463
rect 528944 101453 528954 101463
rect 539544 101460 539554 101470
rect 539934 101460 539944 101470
rect 572544 101463 572554 101473
rect 572934 101463 572944 101473
rect 583544 101463 583554 101473
rect 583934 101463 583944 101473
rect 539534 101450 539544 101460
rect 539944 101450 539954 101460
rect 572534 101453 572544 101463
rect 572944 101453 572954 101463
rect 583534 101453 583544 101463
rect 583944 101453 583954 101463
rect 528534 100962 528544 100972
rect 528944 100962 528954 100972
rect 528544 100952 528554 100962
rect 528934 100952 528944 100962
rect 539534 100961 539544 100971
rect 539944 100961 539954 100971
rect 572534 100962 572544 100972
rect 572944 100962 572954 100972
rect 583534 100962 583544 100972
rect 583944 100962 583954 100972
rect 539544 100951 539554 100961
rect 539934 100951 539944 100961
rect 572544 100952 572554 100962
rect 572934 100952 572944 100962
rect 583544 100952 583554 100962
rect 583934 100952 583944 100962
rect 528544 100591 528554 100601
rect 528934 100591 528944 100601
rect 539544 100597 539554 100607
rect 539934 100597 539944 100607
rect 528534 100581 528544 100591
rect 528944 100581 528954 100591
rect 539534 100587 539544 100597
rect 539944 100587 539954 100597
rect 572544 100596 572554 100606
rect 572934 100596 572944 100606
rect 572534 100586 572544 100596
rect 572944 100586 572954 100596
rect 583544 100595 583554 100605
rect 583934 100595 583944 100605
rect 583534 100585 583544 100595
rect 583944 100585 583954 100595
rect 528534 100026 528544 100036
rect 528944 100026 528954 100036
rect 539534 100029 539544 100039
rect 539944 100029 539954 100039
rect 572534 100029 572544 100039
rect 572944 100029 572954 100039
rect 528544 100016 528554 100026
rect 528934 100016 528944 100026
rect 539544 100019 539554 100029
rect 539934 100019 539944 100029
rect 572544 100019 572554 100029
rect 572934 100019 572944 100029
rect 583534 100027 583544 100037
rect 583944 100027 583954 100037
rect 583544 100017 583554 100027
rect 583934 100017 583944 100027
rect 529284 99648 529294 99658
rect 529674 99648 529684 99658
rect 540284 99648 540294 99658
rect 540674 99648 540684 99658
rect 573284 99648 573294 99658
rect 573674 99648 573684 99658
rect 584284 99648 584294 99658
rect 584674 99648 584684 99658
rect 529274 99638 529284 99648
rect 529684 99638 529694 99648
rect 540274 99638 540284 99648
rect 540684 99638 540694 99648
rect 573274 99638 573284 99648
rect 573684 99638 573694 99648
rect 584274 99638 584284 99648
rect 584684 99638 584694 99648
rect 529274 98726 529284 98736
rect 529684 98726 529694 98736
rect 529284 98716 529294 98726
rect 529674 98716 529684 98726
rect 540274 98725 540284 98735
rect 540684 98725 540694 98735
rect 573274 98731 573284 98741
rect 573684 98731 573694 98741
rect 540284 98715 540294 98725
rect 540674 98715 540684 98725
rect 573284 98721 573294 98731
rect 573674 98721 573684 98731
rect 584274 98726 584284 98736
rect 584684 98726 584694 98736
rect 584284 98716 584294 98726
rect 584674 98716 584684 98726
rect 528544 98259 528554 98269
rect 528934 98259 528944 98269
rect 539544 98265 539554 98275
rect 539934 98265 539944 98275
rect 572544 98265 572554 98275
rect 572934 98265 572944 98275
rect 583544 98265 583554 98275
rect 583934 98265 583944 98275
rect 528534 98249 528544 98259
rect 528944 98249 528954 98259
rect 539534 98255 539544 98265
rect 539944 98255 539954 98265
rect 572534 98255 572544 98265
rect 572944 98255 572954 98265
rect 583534 98255 583544 98265
rect 583944 98255 583954 98265
rect 528534 97305 528544 97315
rect 528944 97305 528954 97315
rect 539534 97311 539544 97321
rect 539944 97311 539954 97321
rect 572534 97311 572544 97321
rect 572944 97311 572954 97321
rect 583534 97312 583544 97322
rect 583944 97312 583954 97322
rect 528544 97295 528554 97305
rect 528934 97295 528944 97305
rect 539544 97301 539554 97311
rect 539934 97301 539944 97311
rect 572544 97301 572554 97311
rect 572934 97301 572944 97311
rect 583544 97302 583554 97312
rect 583934 97302 583944 97312
rect 529284 97094 529294 97104
rect 529674 97094 529684 97104
rect 529274 97084 529284 97094
rect 529684 97084 529694 97094
rect 540284 97087 540294 97097
rect 540674 97087 540684 97097
rect 573284 97091 573294 97101
rect 573674 97091 573684 97101
rect 584284 97091 584294 97101
rect 584674 97091 584684 97101
rect 540274 97077 540284 97087
rect 540684 97077 540694 97087
rect 573274 97081 573284 97091
rect 573684 97081 573694 97091
rect 584274 97081 584284 97091
rect 584684 97081 584694 97091
rect 529274 96730 529284 96740
rect 529684 96730 529694 96740
rect 540274 96730 540284 96740
rect 540684 96730 540694 96740
rect 573274 96730 573284 96740
rect 573684 96730 573694 96740
rect 584274 96730 584284 96740
rect 584684 96730 584694 96740
rect 529284 96720 529294 96730
rect 529674 96720 529684 96730
rect 540284 96720 540294 96730
rect 540674 96720 540684 96730
rect 573284 96720 573294 96730
rect 573674 96720 573684 96730
rect 584284 96720 584294 96730
rect 584674 96720 584684 96730
rect 529284 96263 529294 96273
rect 529674 96263 529684 96273
rect 540284 96263 540294 96273
rect 540674 96263 540684 96273
rect 573284 96263 573294 96273
rect 573674 96263 573684 96273
rect 584284 96263 584294 96273
rect 584674 96263 584684 96273
rect 529274 96253 529284 96263
rect 529684 96253 529694 96263
rect 540274 96253 540284 96263
rect 540684 96253 540694 96263
rect 573274 96253 573284 96263
rect 573684 96253 573694 96263
rect 584274 96253 584284 96263
rect 584684 96253 584694 96263
rect 529274 95960 529284 95970
rect 529684 95960 529694 95970
rect 540274 95960 540284 95970
rect 540684 95960 540694 95970
rect 573274 95960 573284 95970
rect 573684 95960 573694 95970
rect 584274 95961 584284 95971
rect 584684 95961 584694 95971
rect 529284 95950 529294 95960
rect 529674 95950 529684 95960
rect 540284 95950 540294 95960
rect 540674 95950 540684 95960
rect 573284 95950 573294 95960
rect 573674 95950 573684 95960
rect 584284 95951 584294 95961
rect 584674 95951 584684 95961
rect 528544 95869 528554 95879
rect 528934 95869 528944 95879
rect 528534 95859 528544 95869
rect 528944 95859 528954 95869
rect 539544 95864 539554 95874
rect 539934 95864 539944 95874
rect 572544 95864 572554 95874
rect 572934 95864 572944 95874
rect 583544 95868 583554 95878
rect 583934 95868 583944 95878
rect 539534 95854 539544 95864
rect 539944 95854 539954 95864
rect 572534 95854 572544 95864
rect 572944 95854 572954 95864
rect 583534 95858 583544 95868
rect 583944 95858 583954 95868
rect 528534 95551 528544 95561
rect 528944 95551 528954 95561
rect 528544 95541 528554 95551
rect 528934 95541 528944 95551
rect 539534 95545 539544 95555
rect 539944 95545 539954 95555
rect 572534 95549 572544 95559
rect 572944 95549 572954 95559
rect 539544 95535 539554 95545
rect 539934 95535 539944 95545
rect 572544 95539 572554 95549
rect 572934 95539 572944 95549
rect 583534 95547 583544 95557
rect 583944 95547 583954 95557
rect 583544 95537 583554 95547
rect 583934 95537 583944 95547
rect 528544 95156 528554 95166
rect 528934 95156 528944 95166
rect 539544 95162 539554 95172
rect 539934 95162 539944 95172
rect 572544 95162 572554 95172
rect 572934 95162 572944 95172
rect 528534 95146 528544 95156
rect 528944 95146 528954 95156
rect 539534 95152 539544 95162
rect 539944 95152 539954 95162
rect 572534 95152 572544 95162
rect 572944 95152 572954 95162
rect 583544 95161 583554 95171
rect 583934 95161 583944 95171
rect 583534 95151 583544 95161
rect 583944 95151 583954 95161
rect 528534 94841 528544 94851
rect 528944 94841 528954 94851
rect 539534 94843 539544 94853
rect 539944 94843 539954 94853
rect 572534 94843 572544 94853
rect 572944 94843 572954 94853
rect 528544 94831 528554 94841
rect 528934 94831 528944 94841
rect 539544 94833 539554 94843
rect 539934 94833 539944 94843
rect 572544 94833 572554 94843
rect 572934 94833 572944 94843
rect 583534 94842 583544 94852
rect 583944 94842 583954 94852
rect 583544 94832 583554 94842
rect 583934 94832 583944 94842
rect 529284 94642 529294 94652
rect 529674 94642 529684 94652
rect 540284 94642 540294 94652
rect 540674 94642 540684 94652
rect 529274 94632 529284 94642
rect 529684 94632 529694 94642
rect 540274 94632 540284 94642
rect 540684 94632 540694 94642
rect 573284 94640 573294 94650
rect 573674 94640 573684 94650
rect 584284 94640 584294 94650
rect 584674 94640 584684 94650
rect 573274 94630 573284 94640
rect 573684 94630 573694 94640
rect 584274 94630 584284 94640
rect 584684 94630 584694 94640
rect 529274 94396 529284 94406
rect 529684 94396 529694 94406
rect 540274 94398 540284 94408
rect 540684 94398 540694 94408
rect 529284 94386 529294 94396
rect 529674 94386 529684 94396
rect 540284 94388 540294 94398
rect 540674 94388 540684 94398
rect 573274 94394 573284 94404
rect 573684 94394 573694 94404
rect 584274 94396 584284 94406
rect 584684 94396 584694 94406
rect 573284 94384 573294 94394
rect 573674 94384 573684 94394
rect 584284 94386 584294 94396
rect 584674 94386 584684 94396
rect 529284 93999 529294 94009
rect 529674 93999 529684 94009
rect 540284 93999 540294 94009
rect 540674 93999 540684 94009
rect 529274 93989 529284 93999
rect 529684 93989 529694 93999
rect 540274 93989 540284 93999
rect 540684 93989 540694 93999
rect 573284 93998 573294 94008
rect 573674 93998 573684 94008
rect 584284 93998 584294 94008
rect 584674 93998 584684 94008
rect 573274 93988 573284 93998
rect 573684 93988 573694 93998
rect 584274 93988 584284 93998
rect 584684 93988 584694 93998
rect 529274 93748 529284 93758
rect 529684 93748 529694 93758
rect 540274 93748 540284 93758
rect 540684 93748 540694 93758
rect 573274 93748 573284 93758
rect 573684 93748 573694 93758
rect 584274 93748 584284 93758
rect 584684 93748 584694 93758
rect 529284 93738 529294 93748
rect 529674 93738 529684 93748
rect 540284 93738 540294 93748
rect 540674 93738 540684 93748
rect 573284 93738 573294 93748
rect 573674 93738 573684 93748
rect 584284 93738 584294 93748
rect 584674 93738 584684 93748
<< via3 >>
rect 528544 135728 528942 136422
rect 539544 135729 539944 136426
rect 550544 135726 550944 136426
rect 561544 135726 561944 136426
rect 572544 135727 572944 136426
rect 583544 135726 583944 136422
rect 529284 135300 529684 135510
rect 540284 135300 540684 135510
rect 573284 135337 573684 135547
rect 584284 135337 584684 135547
rect 529284 134088 529684 134298
rect 540284 134088 540684 134298
rect 573284 134125 573684 134335
rect 584284 134125 584684 134335
rect 529284 132876 529684 133086
rect 540284 132876 540684 133086
rect 573284 132913 573684 133123
rect 584284 132913 584684 133123
rect 529284 131664 529684 131874
rect 540284 131664 540684 131874
rect 573284 131701 573684 131911
rect 584284 131701 584684 131911
rect 529284 130452 529684 130662
rect 540284 130452 540684 130662
rect 573284 130489 573684 130699
rect 584284 130489 584684 130699
rect 529284 129240 529684 129450
rect 540284 129240 540684 129450
rect 573284 129277 573684 129487
rect 584284 129277 584684 129487
rect 529284 128028 529684 128238
rect 540284 128028 540684 128238
rect 573284 128065 573684 128275
rect 584284 128065 584684 128275
rect 529284 126816 529684 127026
rect 540284 126816 540684 127026
rect 573284 126853 573684 127063
rect 584284 126853 584684 127063
rect 529284 125604 529684 125814
rect 540284 125604 540684 125814
rect 573284 125641 573684 125851
rect 584284 125641 584684 125851
rect 529284 124392 529684 124602
rect 540284 124392 540684 124602
rect 573284 124429 573684 124639
rect 584284 124429 584684 124639
rect 529284 123180 529684 123390
rect 540284 123180 540684 123390
rect 573284 123217 573684 123427
rect 584284 123217 584684 123427
rect 529284 121968 529684 122178
rect 540284 121968 540684 122178
rect 573284 122005 573684 122215
rect 584284 122005 584684 122215
rect 529284 120756 529684 120966
rect 540284 120756 540684 120966
rect 573284 120793 573684 121003
rect 584284 120793 584684 121003
rect 529284 119544 529684 119754
rect 540284 119544 540684 119754
rect 573284 119581 573684 119791
rect 584284 119581 584684 119791
rect 529284 118332 529684 118542
rect 540284 118332 540684 118542
rect 573284 118369 573684 118579
rect 584284 118369 584684 118579
rect 529284 117120 529684 117330
rect 540284 117120 540684 117330
rect 573284 117157 573684 117367
rect 584284 117157 584684 117367
rect 529284 115908 529684 116118
rect 540284 115908 540684 116118
rect 573284 115945 573684 116155
rect 584284 115945 584684 116155
rect 529284 114675 529684 114875
rect 540284 114675 540684 114875
rect 573284 114727 573684 114880
rect 584284 114725 584684 114875
rect 529284 114270 529684 114606
rect 540284 114270 540684 114606
rect 573284 114270 573684 114604
rect 584284 114270 584684 114605
rect 528544 112576 528944 113982
rect 539544 112576 539944 113982
rect 550544 112303 550944 112764
rect 561544 112303 561944 112764
rect 572544 112585 572944 113978
rect 583544 112577 583944 113981
rect 528544 111035 528944 111234
rect 529284 109365 529684 110765
rect 540284 109365 540684 110765
rect 550544 110083 550944 111567
rect 561544 110084 561944 111562
rect 583544 111036 583944 111234
rect 573284 109365 573684 110765
rect 584284 109366 584684 110765
rect 528544 106971 528944 107280
rect 539544 106848 539944 107290
rect 572544 106848 572944 107290
rect 583544 106906 583944 107290
rect 529284 106253 529684 106702
rect 540284 106270 540684 106702
rect 573284 106270 573684 106702
rect 584284 106256 584684 106702
rect 528544 103642 528944 105548
rect 539544 103645 539944 105552
rect 572544 103645 572944 105552
rect 583544 103645 583944 105552
rect 529284 101588 529684 103445
rect 540284 101588 540684 103445
rect 573284 101588 573684 103441
rect 584284 101589 584684 103445
rect 528544 100962 528944 101463
rect 539544 100961 539944 101460
rect 572544 100962 572944 101463
rect 583544 100962 583944 101463
rect 528544 100026 528944 100591
rect 539544 100029 539944 100597
rect 572544 100029 572944 100596
rect 583544 100027 583944 100595
rect 529284 98726 529684 99648
rect 540284 98725 540684 99648
rect 573284 98731 573684 99648
rect 584284 98726 584684 99648
rect 528544 97305 528944 98259
rect 539544 97311 539944 98265
rect 572544 97311 572944 98265
rect 583544 97312 583944 98265
rect 529284 96730 529684 97094
rect 540284 96730 540684 97087
rect 573284 96730 573684 97091
rect 584284 96730 584684 97091
rect 529284 95960 529684 96263
rect 540284 95960 540684 96263
rect 573284 95960 573684 96263
rect 584284 95961 584684 96263
rect 528544 95551 528944 95869
rect 539544 95545 539944 95864
rect 572544 95549 572944 95864
rect 583544 95547 583944 95868
rect 528544 94841 528944 95156
rect 539544 94843 539944 95162
rect 572544 94843 572944 95162
rect 583544 94842 583944 95161
rect 529284 94396 529684 94642
rect 540284 94398 540684 94642
rect 573284 94394 573684 94640
rect 584284 94396 584684 94640
rect 529284 93748 529684 93999
rect 540284 93748 540684 93999
rect 573284 93748 573684 93998
rect 584284 93748 584684 93998
<< end >>
