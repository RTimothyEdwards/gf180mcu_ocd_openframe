magic
tech gf180mcuD
magscale 1 10
timestamp 1765301996
<< checkpaint >>
rect 68239 862158 76146 875981
rect 699782 863562 707769 874986
rect 699762 443741 707799 449816
rect 699935 431181 707819 442391
rect 68178 416034 76187 427409
rect 68128 93100 76186 101937
rect 68210 83087 76268 91924
rect 103118 68166 111952 76196
rect 275710 76169 286982 76248
rect 268113 68150 286982 76169
rect 268113 68139 276947 68150
<< metal4 >>
rect 379272 943800 381172 944000
rect 381752 943800 383802 944000
rect 384122 943800 386172 944000
rect 386828 943800 388878 944000
rect 389198 943800 391248 944000
rect 391828 943800 393728 944000
rect 599272 943800 601172 944000
rect 601752 943800 603802 944000
rect 604122 943800 606172 944000
rect 606828 943800 608878 944000
rect 609198 943800 611248 944000
rect 611828 943800 613728 944000
rect 270272 72147 272172 74169
rect 270272 70567 270282 72147
rect 272162 70567 272172 72147
rect 105272 70000 107172 70200
rect 107752 70000 109802 70200
rect 110122 70000 112172 70200
rect 112828 70000 114878 70200
rect 115198 70000 117248 70200
rect 117828 70000 119728 70200
rect 270272 70000 272172 70567
rect 272752 72147 274802 74169
rect 272752 70567 272762 72147
rect 274792 70567 274802 72147
rect 272752 70000 274802 70567
rect 277828 72147 279878 74248
rect 277828 70567 277838 72147
rect 279868 70567 279878 72147
rect 275122 70000 277172 70200
rect 277828 70000 279878 70567
rect 280198 72147 282248 74248
rect 280198 70567 280208 72147
rect 282238 70567 282248 72147
rect 280198 70000 282248 70567
rect 282828 72147 284728 74248
rect 282828 70567 282838 72147
rect 284718 70567 284728 72147
rect 282828 70000 284728 70567
rect 600272 70000 602172 70200
rect 602752 70000 604802 70200
rect 605122 70000 607172 70200
rect 607828 70000 609878 70200
rect 610198 70000 612248 70200
rect 612828 70000 614728 70200
rect 655272 69999 657172 70199
rect 657752 69999 659802 70199
rect 660122 69999 662172 70199
rect 662828 69999 664878 70199
rect 665198 69999 667248 70199
rect 667828 69999 669728 70199
<< via4 >>
rect 72492 871838 74072 873868
rect 72492 869132 74072 871162
rect 701980 870838 703560 872868
rect 72492 866762 74072 868792
rect 701980 868120 703560 870174
rect 72492 864282 74072 866162
rect 701980 865762 703560 867792
rect 703920 445838 705500 447718
rect 703920 438132 705500 440162
rect 703920 435762 705500 437792
rect 703920 433282 705500 435162
rect 70552 423196 72132 425250
rect 70552 420838 72132 422868
rect 70552 418132 72132 420162
rect 72492 97838 74072 99718
rect 72492 95196 74072 97250
rect 72492 87750 74072 89804
rect 72492 85282 74072 87162
rect 270282 70567 272162 72147
rect 272762 70567 274792 72147
rect 277838 70567 279868 72147
rect 280208 70567 282238 72147
rect 282838 70567 284718 72147
<< metal5 >>
rect 70000 876828 70270 878728
rect 70000 874198 70270 876248
rect 705730 875828 706000 877728
rect 70000 873868 74146 873878
rect 70000 871838 72492 873868
rect 74072 871838 74146 873868
rect 705728 873186 706002 875260
rect 70000 871828 74146 871838
rect 701782 872868 706000 872878
rect 70000 871162 74146 871172
rect 70000 869132 72492 871162
rect 74072 869132 74146 871162
rect 701782 870838 701980 872868
rect 703560 870838 706000 872868
rect 701782 870828 706000 870838
rect 70000 869122 74146 869132
rect 701782 870174 706002 870184
rect 70000 868792 74146 868802
rect 70000 866762 72492 868792
rect 74072 866762 74146 868792
rect 701782 868120 701980 870174
rect 703560 868120 706002 870174
rect 701782 868110 706002 868120
rect 70000 866752 74146 866762
rect 701782 867792 706000 867802
rect 70000 866162 74146 866172
rect 70000 864282 72492 866162
rect 74072 864282 74146 866162
rect 701782 865762 701980 867792
rect 703560 865762 706000 867792
rect 701782 865752 706000 865762
rect 70000 864272 74146 864282
rect 705728 863260 706002 865184
rect 70000 835828 70270 837728
rect 70000 833198 70270 835248
rect 70000 830828 70270 832878
rect 70000 828122 70270 830172
rect 70000 825752 70270 827802
rect 70000 823272 70270 825172
rect 70000 794829 70270 796729
rect 70000 792199 70270 794249
rect 70000 789829 70270 791879
rect 705730 789828 706000 791728
rect 70000 787123 70270 789173
rect 705728 787186 706002 789260
rect 70000 784753 70270 786803
rect 705730 784828 706000 786878
rect 70000 782273 70270 784173
rect 705728 782110 706002 784184
rect 705730 779752 706000 781802
rect 705726 777248 706004 779196
rect 705730 488828 706000 490728
rect 705730 486198 706000 488248
rect 705730 483828 706000 485878
rect 705730 481122 706000 483172
rect 705730 478752 706000 480802
rect 705730 476272 706000 478172
rect 70000 466828 70270 468728
rect 70000 464198 70270 466248
rect 70000 461828 70270 463878
rect 70000 459122 70270 461172
rect 70000 456752 70270 458802
rect 70000 454272 70270 456172
rect 701762 447718 706000 447728
rect 701762 445838 703920 447718
rect 705500 445838 706000 447718
rect 701762 445828 706000 445838
rect 705730 443198 706000 445248
rect 705730 440828 706000 442878
rect 701935 440162 706000 440172
rect 701935 438132 703920 440162
rect 705500 438132 706000 440162
rect 701935 438122 706000 438132
rect 701935 437792 706000 437802
rect 701935 435762 703920 437792
rect 705500 435762 706000 437792
rect 701935 435752 706000 435762
rect 701935 435162 706000 435172
rect 701935 433282 703920 435162
rect 705500 433282 706000 435162
rect 701935 433272 706000 433282
rect 70000 425828 70270 427728
rect 69998 425250 74187 425260
rect 69998 423196 70552 425250
rect 72132 423196 74187 425250
rect 69998 423186 74187 423196
rect 70000 422868 74187 422878
rect 70000 420838 70552 422868
rect 72132 420838 74187 422868
rect 70000 420828 74187 420838
rect 70000 420162 74187 420172
rect 70000 418132 70552 420162
rect 72132 418132 74187 420162
rect 70000 418122 74187 418132
rect 69998 415740 70272 417814
rect 70000 413272 70270 415172
rect 705730 402828 706000 404728
rect 705730 400198 706000 402248
rect 705730 397828 706000 399878
rect 705730 395122 706000 397172
rect 705730 392752 706000 394802
rect 705730 390272 706000 392172
rect 70000 138828 70270 140728
rect 69998 136186 70272 138260
rect 70000 133828 70270 135878
rect 70000 131122 70270 133172
rect 69998 128740 70272 130814
rect 70000 126272 70270 128172
rect 70000 99718 74186 99728
rect 70000 97838 72492 99718
rect 74072 97838 74186 99718
rect 70000 97828 74186 97838
rect 69998 97250 74186 97260
rect 69998 95196 72492 97250
rect 74072 95196 74186 97250
rect 69998 95186 74186 95196
rect 70000 92828 70270 94878
rect 70000 90122 70270 92172
rect 69998 89804 74268 89814
rect 69998 87750 72492 89804
rect 74072 87750 74268 89804
rect 69998 87740 74268 87750
rect 70000 87162 74268 87172
rect 70000 85282 72492 87162
rect 74072 85282 74268 87162
rect 70000 85272 74268 85282
<< comment >>
rect 69593 944007 706407 944407
rect 69593 69993 69993 944007
rect 706007 69993 706407 944007
rect 69593 69593 706407 69993
<< labels >>
flabel metal4 105272 70000 107172 70200 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 107752 70000 109802 70200 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 110122 70000 112172 70200 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 112828 70000 114878 70200 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 115198 70000 117248 70200 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 117828 70000 119728 70200 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 270272 70000 272172 70200 0 FreeSans 1600 0 0 0 vssd
port 625 nsew
flabel metal4 272752 70000 274802 70200 0 FreeSans 1600 0 0 0 vssd
port 625 nsew
flabel metal4 275122 70000 277172 70200 0 FreeSans 1600 0 0 0 vssd
port 625 nsew
flabel metal4 277828 70000 279878 70200 0 FreeSans 1600 0 0 0 vssd
port 625 nsew
flabel metal4 280198 70000 282248 70200 0 FreeSans 1600 0 0 0 vssd
port 625 nsew
flabel metal4 282828 70000 284728 70200 0 FreeSans 1600 0 0 0 vssd
port 625 nsew
flabel metal4 600272 70000 602172 70200 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 602752 70000 604802 70200 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 605122 70000 607172 70200 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 607828 70000 609878 70200 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 610198 70000 612248 70200 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 612828 70000 614728 70200 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 655272 69999 657172 70199 0 FreeSans 1600 0 0 0 vddio
port 626 nsew
flabel metal4 657752 69999 659802 70199 0 FreeSans 1600 0 0 0 vddio
port 626 nsew
flabel metal4 660122 69999 662172 70199 0 FreeSans 1600 0 0 0 vddio
port 626 nsew
flabel metal4 662828 69999 664878 70199 0 FreeSans 1600 0 0 0 vddio
port 626 nsew
flabel metal4 665198 69999 667248 70199 0 FreeSans 1600 0 0 0 vddio
port 626 nsew
flabel metal4 667828 69999 669728 70199 0 FreeSans 1600 0 0 0 vddio
port 626 nsew
flabel metal4 379272 943800 381172 944000 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 381752 943800 383802 944000 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 384122 943800 386172 944000 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 386828 943800 388878 944000 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 389198 943800 391248 944000 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 391828 943800 393728 944000 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 599272 943800 601172 944000 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 601752 943800 603802 944000 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 604122 943800 606172 944000 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 606828 943800 608878 944000 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 609198 943800 611248 944000 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 611828 943800 613728 944000 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal5 705730 390272 706000 392172 0 FreeSans 1600 90 0 0 vssio
port 624 nsew
flabel metal5 705730 392752 706000 394802 0 FreeSans 1600 90 0 0 vssio
port 624 nsew
flabel metal5 705730 395122 706000 397172 0 FreeSans 1600 90 0 0 vssio
port 624 nsew
flabel metal5 705730 397828 706000 399878 0 FreeSans 1600 90 0 0 vssio
port 624 nsew
flabel metal5 705730 400198 706000 402248 0 FreeSans 1600 90 0 0 vssio
port 624 nsew
flabel metal5 705730 402828 706000 404728 0 FreeSans 1600 90 0 0 vssio
port 624 nsew
flabel metal5 705730 433272 706000 435172 0 FreeSans 1600 90 0 0 vssd
port 625 nsew
flabel metal5 705730 435752 706000 437802 0 FreeSans 1600 90 0 0 vssd
port 625 nsew
flabel metal5 705730 438122 706000 440172 0 FreeSans 1600 90 0 0 vssd
port 625 nsew
flabel metal5 705730 440828 706000 442878 0 FreeSans 1600 90 0 0 vssd
port 625 nsew
flabel metal5 705730 443198 706000 445248 0 FreeSans 1600 90 0 0 vssd
port 625 nsew
flabel metal5 705730 445828 706000 447728 0 FreeSans 1600 90 0 0 vssd
port 625 nsew
flabel metal5 705730 476272 706000 478172 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 705730 478752 706000 480802 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 705730 481122 706000 483172 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 705730 483828 706000 485878 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 705730 486198 706000 488248 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 705730 488828 706000 490728 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 705726 777248 706004 779196 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 705730 779752 706000 781802 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 705728 782110 706002 784184 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 705730 784828 706000 786878 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 705728 787186 706002 789260 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 705730 789828 706000 791728 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 705728 863260 706002 865184 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 705730 865752 706000 867802 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 705728 868110 706002 870184 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 705730 870828 706000 872878 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 705728 873186 706002 875260 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 705730 875828 706000 877728 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 70000 85272 70270 87172 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 69998 87740 70272 89814 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 70000 90122 70270 92172 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 70000 92828 70270 94878 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 69998 95186 70272 97260 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 70000 97828 70270 99728 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 70000 126272 70270 128172 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 69998 128740 70272 130814 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 131122 70270 133172 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 133828 70270 135878 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 69998 136186 70272 138260 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 138828 70270 140728 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 413272 70270 415172 0 FreeSans 1600 90 0 0 vssd
port 625 nsew
flabel metal5 69998 415740 70272 417814 0 FreeSans 1600 90 0 0 vssd
port 625 nsew
flabel metal5 70000 418122 70270 420172 0 FreeSans 1600 90 0 0 vssd
port 625 nsew
flabel metal5 70000 420828 70270 422878 0 FreeSans 1600 90 0 0 vssd
port 625 nsew
flabel metal5 69998 423186 70272 425260 0 FreeSans 1600 90 0 0 vssd
port 625 nsew
flabel metal5 70000 425828 70270 427728 0 FreeSans 1600 90 0 0 vssd
port 625 nsew
flabel metal5 70000 454272 70270 456172 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 456752 70270 458802 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 459122 70270 461172 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 461828 70270 463878 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 464198 70270 466248 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 466828 70270 468728 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 782273 70270 784173 0 FreeSans 1600 90 0 0 vssio
port 624 nsew
flabel metal5 70000 784753 70270 786803 0 FreeSans 1600 90 0 0 vssio
port 624 nsew
flabel metal5 70000 787123 70270 789173 0 FreeSans 1600 90 0 0 vssio
port 624 nsew
flabel metal5 70000 789829 70270 791879 0 FreeSans 1600 90 0 0 vssio
port 624 nsew
flabel metal5 70000 792199 70270 794249 0 FreeSans 1600 90 0 0 vssio
port 624 nsew
flabel metal5 70000 794829 70270 796729 0 FreeSans 1600 90 0 0 vssio
port 624 nsew
flabel metal5 70000 823272 70270 825172 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 825752 70270 827802 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 828122 70270 830172 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 830828 70270 832878 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 833198 70270 835248 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 835828 70270 837728 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 864272 70270 866172 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 70000 866752 70270 868802 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 70000 869122 70270 871172 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 70000 871828 70270 873878 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 70000 874198 70270 876248 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 70000 876828 70270 878728 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
<< properties >>
string FIXED_BBOX 70017 70017 705983 943983
<< end >>
