magic
tech gf180mcuD
magscale 1 10
timestamp 1765308861
<< error_p >>
rect -58 -655 -28 -609
<< nwell >>
rect -378 -886 368 886
<< hvpmos >>
rect -60 -576 50 624
<< mvpdiff >>
rect -148 611 -60 624
rect -148 -563 -135 611
rect -89 -563 -60 611
rect -148 -576 -60 -563
rect 50 611 138 624
rect 50 -563 79 611
rect 125 -563 138 611
rect 50 -576 138 -563
<< mvpdiffc >>
rect -135 -563 -89 611
rect 79 -563 125 611
<< mvnsubdiff >>
rect -292 787 282 800
rect -292 741 -169 787
rect 159 741 282 787
rect -292 728 282 741
rect -292 681 -220 728
rect -292 -681 -279 681
rect -233 -681 -220 681
rect 210 681 282 728
rect -292 -728 -220 -681
rect 210 -681 223 681
rect 269 -681 282 681
rect 210 -728 282 -681
rect -292 -800 282 -728
<< mvnsubdiffcont >>
rect -169 741 159 787
rect -279 -681 -233 681
rect 223 -681 269 681
<< polysilicon >>
rect -60 624 50 668
rect -60 -609 50 -576
rect -60 -655 -28 -609
rect 18 -655 50 -609
rect -60 -668 50 -655
<< polycontact >>
rect -28 -655 18 -609
<< metal1 >>
rect -279 741 -169 787
rect 159 741 269 787
rect -279 681 -233 741
rect 223 681 269 741
rect -135 611 -89 622
rect -135 -574 -89 -563
rect 79 611 125 622
rect 79 -574 125 -563
rect -58 -655 -28 -609
rect 18 -655 48 -609
rect -279 -741 -233 -681
rect 223 -741 269 -681
rect -279 -787 269 -741
<< properties >>
string FIXED_BBOX -246 -764 246 764
string GDS_END 38888
string GDS_FILE ../gds/simple_por.gds.gz
string GDS_START 33188
<< end >>
