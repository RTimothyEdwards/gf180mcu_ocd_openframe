magic
tech gf180mcuD
magscale 1 10
timestamp 1765309110
<< metal2 >>
rect 103178 943800 103254 944100
rect 103366 943800 103442 944100
rect 104752 943800 104828 944076
rect 104898 943800 104974 944076
rect 105044 943800 105120 944076
rect 105190 943800 105266 944076
rect 116647 943800 116723 944076
rect 116858 943800 116934 944076
rect 117218 943800 117294 944076
rect 117360 943800 117436 944076
rect 117502 943800 117578 944076
rect 117731 943800 117807 944076
rect 118252 943800 118328 944076
rect 158178 943800 158254 944100
rect 158366 943800 158442 944100
rect 159752 943800 159828 944076
rect 159898 943800 159974 944076
rect 160044 943800 160120 944076
rect 160190 943800 160266 944076
rect 171647 943800 171723 944076
rect 171858 943800 171934 944076
rect 172218 943800 172294 944076
rect 172360 943800 172436 944076
rect 172502 943800 172578 944076
rect 172731 943800 172807 944076
rect 173252 943800 173328 944076
rect 213178 943800 213254 944100
rect 213366 943800 213442 944100
rect 214752 943800 214828 944076
rect 214898 943800 214974 944076
rect 215044 943800 215120 944076
rect 215190 943800 215266 944076
rect 226647 943800 226723 944076
rect 226858 943800 226934 944076
rect 227218 943800 227294 944076
rect 227360 943800 227436 944076
rect 227502 943800 227578 944076
rect 227731 943800 227807 944076
rect 228252 943800 228328 944076
rect 268178 943800 268254 944100
rect 268366 943800 268442 944100
rect 269752 943800 269828 944076
rect 269898 943800 269974 944076
rect 270044 943800 270120 944076
rect 270190 943800 270266 944076
rect 281647 943800 281723 944076
rect 281858 943800 281934 944076
rect 282218 943800 282294 944076
rect 282360 943800 282436 944076
rect 282502 943800 282578 944076
rect 282731 943800 282807 944076
rect 283252 943800 283328 944076
rect 323178 943800 323254 944100
rect 323366 943800 323442 944100
rect 324752 943800 324828 944076
rect 324898 943800 324974 944076
rect 325044 943800 325120 944076
rect 325190 943800 325266 944076
rect 336647 943800 336723 944076
rect 336858 943800 336934 944076
rect 337218 943800 337294 944076
rect 337360 943800 337436 944076
rect 337502 943800 337578 944076
rect 337731 943800 337807 944076
rect 338252 943800 338328 944076
rect 433178 943800 433254 944100
rect 433366 943800 433442 944100
rect 434752 943800 434828 944076
rect 434898 943800 434974 944076
rect 435044 943800 435120 944076
rect 435190 943800 435266 944076
rect 446647 943800 446723 944076
rect 446858 943800 446934 944076
rect 447218 943800 447294 944076
rect 447360 943800 447436 944076
rect 447502 943800 447578 944076
rect 447731 943800 447807 944076
rect 448252 943800 448328 944076
rect 488178 943800 488254 944100
rect 488366 943800 488442 944100
rect 489752 943800 489828 944076
rect 489898 943800 489974 944076
rect 490044 943800 490120 944076
rect 490190 943800 490266 944076
rect 501647 943800 501723 944076
rect 501858 943800 501934 944076
rect 502218 943800 502294 944076
rect 502360 943800 502436 944076
rect 502502 943800 502578 944076
rect 502731 943800 502807 944076
rect 503252 943800 503328 944076
rect 543178 943800 543254 944100
rect 543366 943800 543442 944100
rect 544752 943800 544828 944076
rect 544898 943800 544974 944076
rect 545044 943800 545120 944076
rect 545190 943800 545266 944076
rect 556647 943800 556723 944076
rect 556858 943800 556934 944076
rect 557218 943800 557294 944076
rect 557360 943800 557436 944076
rect 557502 943800 557578 944076
rect 557731 943800 557807 944076
rect 558252 943800 558328 944076
rect 653178 943800 653254 944100
rect 653366 943800 653442 944100
rect 654752 943800 654828 944076
rect 654898 943800 654974 944076
rect 655044 943800 655120 944076
rect 655190 943800 655266 944076
rect 666647 943800 666723 944076
rect 666858 943800 666934 944076
rect 667218 943800 667294 944076
rect 667360 943800 667436 944076
rect 667502 943800 667578 944076
rect 667731 943800 667807 944076
rect 668252 943800 668328 944076
rect 159178 69900 159254 70200
rect 159366 69900 159442 70200
rect 161194 69861 161270 70200
rect 162066 69861 162142 70200
rect 174172 69924 174248 70200
rect 215672 69757 215748 70200
rect 216193 69757 216269 70200
rect 216422 69757 216498 70200
rect 216564 69757 216640 70200
rect 216706 69757 216782 70200
rect 217066 69757 217142 70200
rect 217277 69757 217353 70200
rect 228734 69757 228810 70200
rect 228880 69757 228956 70200
rect 229026 69757 229102 70200
rect 229172 69924 229248 70200
rect 230558 69900 230634 70200
rect 230746 69900 230822 70200
rect 325672 69757 325748 70200
rect 326193 69757 326269 70200
rect 326422 69757 326498 70200
rect 326564 69757 326640 70200
rect 326706 69757 326782 70200
rect 327066 69757 327142 70200
rect 327277 69757 327353 70200
rect 338734 69757 338810 70200
rect 338880 69757 338956 70200
rect 339026 69924 339102 70200
rect 339172 69924 339248 70200
rect 340558 69900 340634 70200
rect 340746 69900 340822 70200
rect 380672 69757 380748 70200
rect 381193 69757 381269 70200
rect 381422 69757 381498 70200
rect 381564 69757 381640 70200
rect 381706 69757 381782 70200
rect 382066 69757 382142 70200
rect 382277 69757 382353 70200
rect 393734 69757 393810 70200
rect 393880 69757 393956 70200
rect 394026 69924 394102 70200
rect 394172 69924 394248 70200
rect 395558 69900 395634 70200
rect 395746 69900 395822 70200
rect 435672 69757 435748 70200
rect 436193 69757 436269 70200
rect 436422 69757 436498 70200
rect 436564 69757 436640 70200
rect 436706 69757 436782 70200
rect 437066 69757 437142 70200
rect 437277 69924 437353 70200
rect 448734 69757 448810 70200
rect 448880 69924 448956 70200
rect 449026 69924 449102 70200
rect 449171 70000 449248 70200
rect 449171 69924 449247 70000
rect 450558 69900 450634 70200
rect 450746 69900 450822 70200
rect 490672 69757 490748 70200
rect 491193 69757 491269 70200
rect 491422 69757 491498 70200
rect 491564 69757 491640 70200
rect 491706 69757 491782 70200
rect 492066 69757 492142 70200
rect 492277 69924 492353 70200
rect 503734 69757 503810 70200
rect 503880 69924 503956 70200
rect 504026 69924 504102 70200
rect 504172 69924 504248 70200
rect 505558 69900 505634 70200
rect 505746 69900 505822 70200
rect 507707 69848 507783 70200
rect 508290 69847 508366 70200
rect 509707 69848 509783 70200
rect 510290 69847 510366 70200
rect 511707 69848 511783 70200
rect 512290 69847 512366 70200
rect 513707 69848 513783 70200
rect 514290 69847 514366 70200
rect 515707 69848 515783 70200
rect 516290 69847 516366 70200
rect 517707 69848 517783 70200
rect 518290 69847 518366 70200
rect 519707 69848 519783 70200
rect 520290 69847 520366 70200
rect 521707 69848 521783 70200
rect 522290 69847 522366 70200
rect 523707 69848 523783 70200
rect 524290 69847 524366 70200
rect 525707 69848 525783 70200
rect 526290 69847 526366 70200
rect 527707 69848 527783 70200
rect 528290 69847 528366 70200
rect 529707 69848 529783 70200
rect 530290 69847 530366 70200
rect 531707 69848 531783 70200
rect 532290 69847 532366 70200
rect 533707 69848 533783 70200
rect 534290 69847 534366 70200
rect 535707 69848 535783 70200
rect 536290 69847 536366 70200
rect 537707 69848 537783 70200
rect 538290 69847 538366 70200
rect 545672 69924 545748 70200
rect 546193 69924 546269 70200
rect 546422 69924 546498 70200
rect 546564 69923 546640 70200
rect 546706 69923 546782 70200
rect 547066 69924 547142 70200
rect 547277 69924 547353 70200
rect 558734 69924 558810 70200
rect 558880 69924 558956 70200
rect 559026 69924 559102 70200
rect 559172 69924 559248 70200
rect 560558 69900 560634 70200
rect 560746 69900 560822 70200
rect 590707 69839 590783 70200
rect 590707 69721 590763 69839
rect 591290 69762 591366 70200
rect 593218 69829 593294 70200
rect 591290 69706 592715 69762
rect 507707 9592 507763 13172
rect 508290 9704 508346 13172
rect 509707 9816 509763 13172
rect 510290 9928 510346 13172
rect 511707 10041 511763 13172
rect 512290 10153 512346 13172
rect 512717 12684 512918 13624
rect 512717 11773 512729 12684
rect 512898 11773 512918 12684
rect 512717 11751 512918 11773
rect 513081 12684 513282 13624
rect 513081 11773 513095 12684
rect 513264 11773 513282 12684
rect 513081 11751 513282 11773
rect 513707 10265 513763 13172
rect 514290 10377 514346 13172
rect 515707 10489 515763 13172
rect 516290 10601 516346 13172
rect 517707 10713 517763 13172
rect 517860 12685 518211 14292
rect 517860 11772 517876 12685
rect 518165 11772 518211 12685
rect 517860 11751 518211 11772
rect 518290 10825 518346 13172
rect 519707 10825 519763 13172
rect 520290 10825 520346 13172
rect 521707 10825 521763 13172
rect 522290 10825 522346 13172
rect 522717 12685 522918 13642
rect 522717 11772 522731 12685
rect 522905 11772 522918 12685
rect 522717 11751 522918 11772
rect 523081 12686 523282 13642
rect 523081 11773 523097 12686
rect 523271 11773 523282 12686
rect 523081 11751 523282 11773
rect 523707 11273 523763 13172
rect 518290 10769 519466 10825
rect 519707 10769 520138 10825
rect 520290 10769 520810 10825
rect 517707 10657 518682 10713
rect 516290 10545 518010 10601
rect 515707 10488 517309 10489
rect 515707 10433 517338 10488
rect 514290 10321 516666 10377
rect 513707 10209 515882 10265
rect 512290 10097 515210 10153
rect 511707 9985 514538 10041
rect 510290 9872 513866 9928
rect 509707 9760 513194 9816
rect 508290 9648 512410 9704
rect 507707 9536 511738 9592
rect 512354 9518 512410 9648
rect 513138 9504 513194 9760
rect 513810 9535 513866 9872
rect 514482 9536 514538 9985
rect 515154 9536 515210 10097
rect 515826 9536 515882 10209
rect 516610 9531 516666 10321
rect 517282 9528 517338 10433
rect 517954 9536 518010 10545
rect 518626 9536 518682 10657
rect 519410 9535 519466 10769
rect 520082 9536 520138 10769
rect 520754 9528 520810 10769
rect 521426 10769 521763 10825
rect 522098 10769 522346 10825
rect 522882 11217 523763 11273
rect 521426 9502 521482 10769
rect 522098 9536 522154 10769
rect 522882 9536 522938 11217
rect 524290 11161 524346 13172
rect 523554 11105 524346 11161
rect 523554 9536 523610 11105
rect 525707 11049 525763 13172
rect 525860 12942 526211 14305
rect 525860 11780 525881 12942
rect 526166 11780 526211 12942
rect 525860 11751 526211 11780
rect 524226 10993 525763 11049
rect 524226 9536 524282 10993
rect 526290 10937 526346 13172
rect 524898 10881 526346 10937
rect 524898 9536 524954 10881
rect 527707 10825 527763 13172
rect 525682 10769 527763 10825
rect 525682 9536 525738 10769
rect 528290 10713 528346 13172
rect 526354 10657 528346 10713
rect 526354 9536 526410 10657
rect 529707 10601 529763 13172
rect 527026 10545 529763 10601
rect 527026 9536 527082 10545
rect 530290 10489 530346 13172
rect 530717 12692 530918 13662
rect 530717 11736 530728 12692
rect 530900 11736 530918 12692
rect 530717 11689 530918 11736
rect 531081 12694 531282 13662
rect 531081 11738 531093 12694
rect 531265 11738 531282 12694
rect 531081 11689 531282 11738
rect 527698 10433 530346 10489
rect 527698 9536 527754 10433
rect 531707 10377 531763 13172
rect 528370 10321 531763 10377
rect 528370 9536 528426 10321
rect 532290 10265 532346 13172
rect 529154 10209 532346 10265
rect 529154 9536 529210 10209
rect 533707 10153 533763 13172
rect 529826 10097 533763 10153
rect 529826 9536 529882 10097
rect 534290 10041 534346 13172
rect 530498 9985 534346 10041
rect 530498 9536 530554 9985
rect 535707 9928 535763 13172
rect 531170 9872 535763 9928
rect 531170 9536 531226 9872
rect 536290 9816 536346 13172
rect 531954 9760 536346 9816
rect 531954 9536 532010 9760
rect 537707 9704 537763 13172
rect 532626 9648 537763 9704
rect 532626 9536 532682 9648
rect 538290 9592 538346 13172
rect 568418 9752 568694 23581
rect 569349 11533 569591 14049
rect 569250 11480 570030 11533
rect 569250 10827 569304 11480
rect 569986 10827 570030 11480
rect 569250 10775 570030 10827
rect 570418 9752 570694 23581
rect 571349 11535 571591 14049
rect 571108 11480 571888 11535
rect 571108 10827 571167 11480
rect 571849 10827 571888 11480
rect 571108 10777 571888 10827
rect 572418 9752 572694 23581
rect 573349 11535 573591 14049
rect 573096 11476 573876 11535
rect 573096 10823 573149 11476
rect 573831 10823 573876 11476
rect 573096 10777 573876 10823
rect 574418 9752 574694 23581
rect 575349 11535 575591 14049
rect 575002 11483 575778 11535
rect 575002 10830 575049 11483
rect 575731 10830 575778 11483
rect 575002 10777 575778 10830
rect 590707 10506 590763 13403
rect 591290 10659 591346 13368
rect 591290 10603 592837 10659
rect 590707 10450 592705 10506
rect 533298 9536 538346 9592
rect 568414 9168 574697 9752
rect 568414 9167 570164 9168
rect 570753 9167 574697 9168
rect 592649 8173 592705 10450
rect 592113 8117 592705 8173
rect 592781 7728 592837 10603
rect 592099 7672 592837 7728
<< via2 >>
rect 512729 11773 512898 12684
rect 513095 11773 513264 12684
rect 517876 11772 518165 12685
rect 522731 11772 522905 12685
rect 523097 11773 523271 12686
rect 525881 11780 526166 12942
rect 530728 11736 530900 12692
rect 531093 11738 531265 12694
rect 569304 10827 569986 11480
rect 571167 10827 571849 11480
rect 573149 10823 573831 11476
rect 575049 10830 575731 11483
<< metal3 >>
rect 705729 921746 706029 921822
rect 705729 921558 706029 921634
rect 705729 920172 706005 920248
rect 705729 920026 706005 920102
rect 705729 919880 706005 919956
rect 705729 919734 706005 919810
rect 69995 919252 70271 919328
rect 69995 918731 70271 918807
rect 69995 918502 70271 918578
rect 69995 918360 70271 918436
rect 69995 918218 70271 918294
rect 69995 917858 70271 917934
rect 69995 917647 70271 917723
rect 705729 908277 706005 908353
rect 705729 908066 706005 908142
rect 705729 907706 706005 907782
rect 705729 907564 706005 907640
rect 705729 907422 706005 907498
rect 705729 907193 706005 907269
rect 705729 906672 706005 906748
rect 69995 906190 70271 906266
rect 69995 906044 70271 906120
rect 69995 905898 70271 905974
rect 69995 905752 70271 905828
rect 69971 904366 70271 904442
rect 69971 904178 70271 904254
rect 705729 835746 706029 835822
rect 705729 835558 706029 835634
rect 705729 834172 706005 834248
rect 705729 834026 706005 834102
rect 705729 833880 706005 833956
rect 705729 833734 706005 833810
rect 705729 822277 706005 822353
rect 705729 822066 706005 822142
rect 705729 821706 706005 821782
rect 705729 821564 706005 821640
rect 705729 821422 706005 821498
rect 705729 821193 706005 821269
rect 705729 820672 706005 820748
rect 69995 755252 70271 755328
rect 69995 754731 70271 754807
rect 69995 754502 70271 754578
rect 69995 754360 70271 754436
rect 69995 754218 70271 754294
rect 69995 753858 70271 753934
rect 69995 753647 70271 753723
rect 705729 749746 706029 749822
rect 705729 749558 706029 749634
rect 705729 748172 706005 748248
rect 705729 748026 706005 748102
rect 705729 747880 706005 747956
rect 705729 747734 706005 747810
rect 69995 742190 70271 742266
rect 69995 742044 70271 742120
rect 69995 741898 70271 741974
rect 69995 741752 70271 741828
rect 69971 740366 70271 740442
rect 69971 740178 70271 740254
rect 705729 736277 706005 736353
rect 705729 736066 706005 736142
rect 705729 735706 706005 735782
rect 705729 735564 706005 735640
rect 705729 735422 706005 735498
rect 705729 735193 706005 735269
rect 705729 734672 706005 734748
rect 69995 714252 70271 714328
rect 69995 713731 70271 713807
rect 69995 713502 70271 713578
rect 69995 713360 70271 713436
rect 69995 713218 70271 713294
rect 69995 712858 70271 712934
rect 69995 712647 70271 712723
rect 705729 706746 706029 706822
rect 705729 706558 706029 706634
rect 705729 705172 706005 705248
rect 705729 705026 706005 705102
rect 705729 704880 706005 704956
rect 705729 704734 706005 704810
rect 69995 701190 70271 701266
rect 69995 701044 70271 701120
rect 69995 700898 70271 700974
rect 69995 700752 70271 700828
rect 69971 699366 70271 699442
rect 69971 699178 70271 699254
rect 705729 693277 706005 693353
rect 705729 693066 706005 693142
rect 705729 692706 706005 692782
rect 705729 692564 706005 692640
rect 705729 692422 706005 692498
rect 705729 692193 706005 692269
rect 705729 691672 706005 691748
rect 69995 673252 70271 673328
rect 69995 672731 70271 672807
rect 69995 672502 70271 672578
rect 69995 672360 70271 672436
rect 69995 672218 70271 672294
rect 69995 671858 70271 671934
rect 69995 671647 70271 671723
rect 705729 663746 706029 663822
rect 705729 663558 706029 663634
rect 705729 662172 706005 662248
rect 705729 662026 706005 662102
rect 705729 661880 706005 661956
rect 705729 661734 706005 661810
rect 69995 660190 70271 660266
rect 69995 660044 70271 660120
rect 69995 659898 70271 659974
rect 69995 659752 70271 659828
rect 69971 658366 70271 658442
rect 69971 658178 70271 658254
rect 705729 650277 706005 650353
rect 705729 650066 706005 650142
rect 705729 649706 706005 649782
rect 705729 649564 706005 649640
rect 705729 649422 706005 649498
rect 705729 649193 706005 649269
rect 705729 648672 706005 648748
rect 69995 632252 70271 632328
rect 69995 631731 70271 631807
rect 69995 631502 70271 631578
rect 69995 631360 70271 631436
rect 69995 631218 70271 631294
rect 69995 630858 70271 630934
rect 69995 630647 70271 630723
rect 705729 620746 706029 620822
rect 705729 620558 706029 620634
rect 69995 619190 70271 619266
rect 705729 619172 706005 619248
rect 69995 619044 70271 619120
rect 705729 619026 706005 619102
rect 69995 618898 70271 618974
rect 705729 618880 706005 618956
rect 69995 618752 70271 618828
rect 705729 618734 706005 618810
rect 69971 617366 70271 617442
rect 69971 617178 70271 617254
rect 705729 607277 706005 607353
rect 705729 607066 706005 607142
rect 705729 606706 706005 606782
rect 705729 606564 706005 606640
rect 705729 606422 706005 606498
rect 705729 606193 706005 606269
rect 705729 605672 706005 605748
rect 69995 591252 70271 591328
rect 69995 590731 70271 590807
rect 69995 590502 70271 590578
rect 69995 590360 70271 590436
rect 69995 590218 70271 590294
rect 69995 589858 70271 589934
rect 69995 589647 70271 589723
rect 69995 578190 70271 578266
rect 69995 578044 70271 578120
rect 69995 577898 70271 577974
rect 69995 577752 70271 577828
rect 705729 577746 706029 577822
rect 705729 577558 706029 577634
rect 69971 576366 70271 576442
rect 69971 576178 70271 576254
rect 705729 576172 706005 576248
rect 705729 576026 706005 576102
rect 705729 575880 706005 575956
rect 705729 575734 706005 575810
rect 705729 564277 706005 564353
rect 705729 564066 706005 564142
rect 705729 563706 706005 563782
rect 705729 563564 706005 563640
rect 705729 563422 706005 563498
rect 705729 563193 706005 563269
rect 705729 562672 706005 562748
rect 69995 550252 70271 550328
rect 69995 549731 70271 549807
rect 69995 549502 70271 549578
rect 69995 549360 70271 549436
rect 69995 549218 70271 549294
rect 69995 548858 70271 548934
rect 69995 548647 70271 548723
rect 69995 537190 70271 537266
rect 69995 537044 70271 537120
rect 69995 536898 70271 536974
rect 69995 536752 70271 536828
rect 69971 535366 70271 535442
rect 69971 535178 70271 535254
rect 705729 534746 706029 534822
rect 705729 534558 706029 534634
rect 705729 533172 706005 533248
rect 705729 533026 706005 533102
rect 705729 532880 706005 532956
rect 705729 532734 706005 532810
rect 705729 521277 706005 521353
rect 705729 521066 706005 521142
rect 705729 520706 706005 520782
rect 705729 520564 706005 520640
rect 705729 520422 706005 520498
rect 705729 520193 706005 520269
rect 705729 519672 706005 519748
rect 69995 509252 70271 509328
rect 69995 508731 70271 508807
rect 69995 508502 70271 508578
rect 69995 508360 70271 508436
rect 69995 508218 70271 508294
rect 69995 507858 70271 507934
rect 69995 507647 70271 507723
rect 69995 496190 70271 496266
rect 69995 496044 70271 496120
rect 69995 495898 70271 495974
rect 69995 495752 70271 495828
rect 69971 494366 70271 494442
rect 69971 494178 70271 494254
rect 69995 386252 70271 386328
rect 69995 385731 70271 385807
rect 69995 385502 70271 385578
rect 69995 385360 70271 385436
rect 69995 385218 70271 385294
rect 69995 384858 70271 384934
rect 69995 384647 70271 384723
rect 69995 373190 70271 373266
rect 69995 373044 70271 373120
rect 69995 372898 70271 372974
rect 69995 372752 70271 372828
rect 69971 371366 70271 371442
rect 69971 371178 70271 371254
rect 705729 362746 706029 362822
rect 705729 362558 706029 362634
rect 705729 361172 706005 361248
rect 705729 361026 706005 361102
rect 705729 360880 706005 360956
rect 705729 360734 706005 360810
rect 705729 349277 706005 349353
rect 705729 349066 706005 349142
rect 705729 348706 706005 348782
rect 705729 348564 706005 348640
rect 705729 348422 706005 348498
rect 705729 348193 706005 348269
rect 705729 347672 706005 347748
rect 69995 345252 70271 345328
rect 69995 344731 70271 344807
rect 69995 344502 70271 344578
rect 69995 344360 70271 344436
rect 69995 344218 70271 344294
rect 69995 343858 70271 343934
rect 69995 343647 70271 343723
rect 69995 332190 70271 332266
rect 69995 332044 70271 332120
rect 69995 331898 70271 331974
rect 69995 331752 70271 331828
rect 69971 330366 70271 330442
rect 69971 330178 70271 330254
rect 705729 319746 706029 319822
rect 705729 319558 706029 319634
rect 705729 318172 706005 318248
rect 705729 318026 706005 318102
rect 705729 317880 706005 317956
rect 705729 317734 706005 317810
rect 705729 306277 706005 306353
rect 705729 306066 706005 306142
rect 705729 305706 706005 305782
rect 705729 305564 706005 305640
rect 705729 305422 706005 305498
rect 705729 305193 706005 305269
rect 705729 304672 706005 304748
rect 69995 304252 70271 304328
rect 69995 303731 70271 303807
rect 69995 303502 70271 303578
rect 69995 303360 70271 303436
rect 69995 303218 70271 303294
rect 69995 302858 70271 302934
rect 69995 302647 70271 302723
rect 69995 291190 70271 291266
rect 69995 291044 70271 291120
rect 69995 290898 70271 290974
rect 69995 290752 70271 290828
rect 69971 289366 70271 289442
rect 69971 289178 70271 289254
rect 705729 276746 706029 276822
rect 705729 276558 706029 276634
rect 705729 275172 706005 275248
rect 705729 275026 706005 275102
rect 705729 274880 706005 274956
rect 705729 274734 706005 274810
rect 69995 263252 70271 263328
rect 705729 263277 706005 263353
rect 705729 263066 706005 263142
rect 69995 262731 70271 262807
rect 705729 262706 706005 262782
rect 69995 262502 70271 262578
rect 705729 262564 706005 262640
rect 69995 262360 70271 262436
rect 705729 262422 706005 262498
rect 69995 262218 70271 262294
rect 705729 262193 706005 262269
rect 69995 261858 70271 261934
rect 69995 261647 70271 261723
rect 705729 261672 706005 261748
rect 69995 250190 70271 250266
rect 69995 250044 70271 250120
rect 69995 249898 70271 249974
rect 69995 249752 70271 249828
rect 69971 248366 70271 248442
rect 69971 248178 70271 248254
rect 705729 233746 706029 233822
rect 705729 233558 706029 233634
rect 705729 232172 706005 232248
rect 705729 232026 706005 232102
rect 705729 231880 706005 231956
rect 705729 231734 706005 231810
rect 69995 222252 70271 222328
rect 69995 221731 70271 221807
rect 69995 221502 70271 221578
rect 69995 221360 70271 221436
rect 69995 221218 70271 221294
rect 69995 220858 70271 220934
rect 69995 220647 70271 220723
rect 705729 220277 706005 220353
rect 705729 220066 706005 220142
rect 705729 219706 706005 219782
rect 705729 219564 706005 219640
rect 705729 219422 706005 219498
rect 705729 219193 706005 219269
rect 705729 218672 706005 218748
rect 69995 209190 70271 209266
rect 69995 209044 70271 209120
rect 69995 208898 70271 208974
rect 69995 208752 70271 208828
rect 69971 207366 70271 207442
rect 69971 207178 70271 207254
rect 705729 190746 706029 190822
rect 705729 190558 706029 190634
rect 705729 189172 706005 189248
rect 705729 189026 706005 189102
rect 705729 188880 706005 188956
rect 705729 188734 706005 188810
rect 69995 181252 70271 181328
rect 69995 180731 70271 180807
rect 69995 180502 70271 180578
rect 69995 180360 70271 180436
rect 69995 180218 70271 180294
rect 69995 179858 70271 179934
rect 69995 179647 70271 179723
rect 705729 177277 706005 177353
rect 705729 177066 706005 177142
rect 705729 176706 706005 176782
rect 705729 176564 706005 176640
rect 705729 176422 706005 176498
rect 705729 176193 706005 176269
rect 705729 175672 706005 175748
rect 69995 168190 70271 168266
rect 69995 168044 70271 168120
rect 69995 167898 70271 167974
rect 69995 167752 70271 167828
rect 69971 166366 70271 166442
rect 69971 166178 70271 166254
rect 705729 147746 706029 147822
rect 705729 147558 706029 147634
rect 705730 146172 706119 146248
rect 705730 146026 706119 146102
rect 705730 145880 706119 145956
rect 705730 145734 706119 145810
rect 705729 134277 706128 134353
rect 705729 134066 706128 134142
rect 705729 133706 706107 133782
rect 705729 133564 706128 133640
rect 705729 133422 706128 133498
rect 705729 133193 706128 133269
rect 705729 132672 706128 132748
rect 705729 104746 706029 104822
rect 705729 104558 706029 104634
rect 705729 103172 706005 103248
rect 705729 103026 706005 103102
rect 705729 102880 706005 102956
rect 705729 102734 706005 102810
rect 705729 91277 706005 91353
rect 705729 91066 706005 91142
rect 705729 90706 706005 90782
rect 705729 90564 706005 90640
rect 705729 90422 706005 90498
rect 705729 90193 706005 90269
rect 705729 89672 706005 89748
rect 525862 12942 526192 12957
rect 512715 12684 513280 12707
rect 512715 11773 512729 12684
rect 512898 11773 513095 12684
rect 513264 11773 513280 12684
rect 512715 11753 513280 11773
rect 517851 12685 518181 12703
rect 517851 11772 517876 12685
rect 518165 11772 518181 12685
rect 512847 10933 513177 11753
rect 512847 10603 513681 10933
rect 513351 9338 513681 10603
rect 517851 9338 518181 11772
rect 522411 12702 522741 12703
rect 522411 12686 523282 12702
rect 522411 12685 523097 12686
rect 522411 11772 522731 12685
rect 522905 11773 523097 12685
rect 523271 11773 523282 12686
rect 522905 11772 523282 11773
rect 522411 11753 523282 11772
rect 525862 11780 525881 12942
rect 526166 11780 526192 12942
rect 522411 9338 522741 11753
rect 525862 11439 526192 11780
rect 530720 12703 531469 12704
rect 530720 12694 531661 12703
rect 530720 12692 531093 12694
rect 530720 11736 530728 12692
rect 530900 11738 531093 12692
rect 531265 11738 531661 12694
rect 530900 11736 531661 11738
rect 530720 11722 531661 11736
rect 525862 11109 527181 11439
rect 526851 9338 527181 11109
rect 531331 9338 531661 11722
rect 569251 11498 575779 11534
rect 569251 10821 569296 11498
rect 569955 11483 575779 11498
rect 569955 11480 575049 11483
rect 569986 10827 571167 11480
rect 571849 11476 575049 11480
rect 571849 10827 573149 11476
rect 569955 10823 573149 10827
rect 573831 10830 575049 11476
rect 575731 10830 575779 11483
rect 573831 10823 575779 10830
rect 569955 10821 575779 10823
rect 569251 10776 575779 10821
<< via3 >>
rect 569296 11480 569955 11498
rect 569296 10827 569304 11480
rect 569304 10827 569955 11480
rect 569296 10821 569955 10827
<< metal4 >>
rect 379272 943800 381172 944000
rect 381752 943800 383802 944000
rect 384122 943800 386172 944000
rect 386828 943800 388878 944000
rect 389198 943800 391248 944000
rect 391828 943800 393728 944000
rect 599272 943800 601172 944000
rect 601752 943800 603802 944000
rect 604122 943800 606172 944000
rect 606828 943800 608878 944000
rect 609198 943800 611248 944000
rect 611828 943800 613728 944000
rect 105272 70000 107172 70200
rect 107752 70000 109802 70200
rect 110122 70000 112172 70200
rect 112828 70000 114878 70200
rect 115198 70000 117248 70200
rect 117828 70000 119728 70200
rect 270272 70000 272172 70200
rect 272752 70000 274802 70200
rect 275122 70000 277172 70200
rect 277828 70000 279878 70200
rect 280198 70000 282248 70200
rect 282828 70000 284728 70200
rect 600272 70000 602172 70200
rect 602752 70000 604802 70200
rect 605122 70000 607172 70200
rect 607828 70000 609878 70200
rect 610198 70000 612248 70200
rect 612828 70000 614728 70200
rect 655272 69999 657172 70199
rect 657752 69999 659802 70199
rect 660122 69999 662172 70199
rect 662828 69999 664878 70199
rect 665198 69999 667248 70199
rect 667828 69999 669728 70199
rect 569251 11498 570004 11529
rect 569251 10821 569296 11498
rect 569955 10821 570004 11498
rect 569251 7878 570004 10821
rect 569251 7125 571348 7878
<< metal5 >>
rect 105500 1001600 117500 1013600
rect 160500 1001600 172500 1013600
rect 215500 1001600 227500 1013600
rect 270500 1001600 282500 1013600
rect 325500 1001600 337500 1013600
rect 380500 1001600 392500 1013600
rect 435500 1001600 447500 1013600
rect 490500 1001600 502500 1013600
rect 545500 1001600 557500 1013600
rect 600500 1001600 612500 1013600
rect 655500 1001600 667500 1013600
rect 400 906500 12400 918500
rect 763600 907500 775600 919500
rect 400 865500 12400 877500
rect 70000 876828 70271 878728
rect 70000 874198 70271 876248
rect 705730 875828 706000 877728
rect 70000 871828 70271 873878
rect 705730 873198 706000 875248
rect 70000 869122 70271 871172
rect 705730 870828 706000 872878
rect 70000 866752 70271 868802
rect 705730 868122 706000 870172
rect 70000 864272 70271 866172
rect 705730 865752 706000 867802
rect 705730 863272 706000 865172
rect 763600 864500 775600 876500
rect 400 824500 12400 836500
rect 70000 835828 70270 837728
rect 70000 833198 70270 835248
rect 70000 830828 70270 832878
rect 70000 828122 70270 830172
rect 70000 825752 70270 827802
rect 70000 823272 70270 825172
rect 763600 821500 775600 833500
rect 400 783500 12400 795500
rect 70000 794829 70270 796729
rect 70000 792199 70270 794249
rect 70000 789829 70270 791879
rect 705730 789828 706000 791728
rect 70000 787123 70270 789173
rect 705730 787198 706000 789248
rect 70000 784753 70270 786803
rect 705730 784828 706000 786878
rect 70000 782273 70270 784173
rect 705730 782122 706000 784172
rect 705730 779752 706000 781802
rect 705730 777272 706000 779172
rect 763600 778500 775600 790500
rect 400 742500 12400 754500
rect 763600 735500 775600 747500
rect 400 701500 12400 713500
rect 763600 692500 775600 704500
rect 400 660500 12400 672500
rect 763600 649500 775600 661500
rect 400 619500 12400 631500
rect 763600 606500 775600 618500
rect 400 578500 12400 590500
rect 763600 563500 775600 575500
rect 400 537500 12400 549500
rect 763600 520500 775600 532500
rect 400 496500 12400 508500
rect 705730 488828 706000 490728
rect 705730 486198 706000 488248
rect 705730 483828 706000 485878
rect 705730 481122 706000 483172
rect 705730 478752 706000 480802
rect 705730 476272 706000 478172
rect 763600 477500 775600 489500
rect 400 455500 12400 467500
rect 70000 466828 70270 468728
rect 70000 464198 70270 466248
rect 70000 461828 70270 463878
rect 70000 459122 70270 461172
rect 70000 456752 70270 458802
rect 70000 454272 70270 456172
rect 705730 445828 706000 447728
rect 705730 443198 706000 445248
rect 705730 440828 706000 442878
rect 705730 438122 706000 440172
rect 705730 435752 706000 437802
rect 705730 433272 706000 435172
rect 763600 434500 775600 446500
rect 400 414500 12400 426500
rect 70000 425828 70270 427728
rect 70000 423198 70270 425248
rect 70000 420828 70270 422878
rect 70000 418122 70270 420172
rect 70000 415752 70270 417802
rect 70000 413272 70270 415172
rect 705730 402828 706000 404728
rect 705730 400198 706000 402248
rect 705730 397828 706000 399878
rect 705730 395122 706000 397172
rect 705730 392752 706000 394802
rect 705730 390272 706000 392172
rect 763600 391500 775600 403500
rect 400 373500 12400 385500
rect 763600 348500 775600 360500
rect 400 332500 12400 344500
rect 763600 305500 775600 317500
rect 400 291500 12400 303500
rect 763600 262500 775600 274500
rect 400 250500 12400 262500
rect 400 209500 12400 221500
rect 763600 219500 775600 231500
rect 400 168500 12400 180500
rect 763600 176500 775600 188500
rect 400 127500 12400 139500
rect 70000 138828 70270 140728
rect 70000 136198 70270 138248
rect 70000 133828 70270 135878
rect 763600 133500 775600 145500
rect 70000 131122 70270 133172
rect 70000 128752 70270 130802
rect 70000 126272 70270 128172
rect 400 86500 12400 98500
rect 70000 97828 70270 99728
rect 70000 95198 70270 97248
rect 70000 92828 70270 94878
rect 70000 90122 70270 92172
rect 763600 90500 775600 102500
rect 70000 87752 70270 89802
rect 70000 85272 70270 87172
rect 106500 400 118500 12400
rect 161500 400 173500 12400
rect 216500 400 228500 12400
rect 271500 400 283500 12400
rect 326500 400 338500 12400
rect 381500 400 393500 12400
rect 436500 400 448500 12400
rect 491500 400 503500 12400
rect 546500 400 558500 12400
rect 601500 400 613500 12400
rect 656500 400 668500 12400
<< comment >>
rect 70013 943983 705987 943987
rect 70013 70017 70017 943983
rect 705983 70017 705987 943983
rect 70013 70013 175579 70017
rect 175817 70013 705987 70017
use gf180mcu_ocd_io__cor  corner[0] $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765222618
transform 1 0 0 0 1 0
box 13097 13097 71000 71000
use gf180mcu_ocd_io__cor  corner[1]
timestamp 1765222618
transform -1 0 776000 0 1 0
box 13097 13097 71000 71000
use gf180mcu_ocd_io__bi_a  gf180mcu_ocd_io__bi_a_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765222618
transform 1 0 215000 0 1 0
box -32 0 15032 70001
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765222618
transform 1 0 704000 0 1 0
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_1
timestamp 1765222618
transform -1 0 72000 0 -1 1014000
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill5  gf180mcu_ocd_io__fill5_2
timestamp 1765222618
transform 0 1 0 -1 0 943000
box -32 13097 1032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765222618
transform 1 0 175000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1
timestamp 1765222618
transform 1 0 71000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_2
timestamp 1765222618
transform 1 0 73000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_3
timestamp 1765222618
transform 1 0 75000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_4
timestamp 1765222618
transform 1 0 77000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_5
timestamp 1765222618
transform 1 0 79000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_6
timestamp 1765222618
transform 1 0 81000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_7
timestamp 1765222618
transform 1 0 83000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_8
timestamp 1765222618
transform 1 0 85000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_9
timestamp 1765222618
transform 1 0 87000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_10
timestamp 1765222618
transform 1 0 89000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_11
timestamp 1765222618
transform 1 0 91000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_12
timestamp 1765222618
transform 1 0 93000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_13
timestamp 1765222618
transform 1 0 95000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_14
timestamp 1765222618
transform 1 0 97000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_15
timestamp 1765222618
transform 1 0 99000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_16
timestamp 1765222618
transform 1 0 101000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_17
timestamp 1765222618
transform 1 0 103000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_18
timestamp 1765222618
transform 1 0 120000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_19
timestamp 1765222618
transform 1 0 122000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_20
timestamp 1765222618
transform 1 0 124000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_21
timestamp 1765222618
transform 1 0 126000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_22
timestamp 1765222618
transform 1 0 128000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_23
timestamp 1765222618
transform 1 0 130000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_24
timestamp 1765222618
transform 1 0 132000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_25
timestamp 1765222618
transform 1 0 134000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_26
timestamp 1765222618
transform 1 0 136000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_27
timestamp 1765222618
transform 1 0 138000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_28
timestamp 1765222618
transform 1 0 140000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_29
timestamp 1765222618
transform 1 0 142000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_30
timestamp 1765222618
transform 1 0 144000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_31
timestamp 1765222618
transform 1 0 146000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_32
timestamp 1765222618
transform 1 0 148000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_33
timestamp 1765222618
transform 1 0 150000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_34
timestamp 1765222618
transform 1 0 152000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_35
timestamp 1765222618
transform 1 0 154000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_36
timestamp 1765222618
transform 1 0 156000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_39
timestamp 1765222618
transform 1 0 177000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_40
timestamp 1765222618
transform 1 0 179000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_41
timestamp 1765222618
transform 1 0 181000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_42
timestamp 1765222618
transform 1 0 183000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_43
timestamp 1765222618
transform 1 0 185000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_44
timestamp 1765222618
transform 1 0 187000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_45
timestamp 1765222618
transform 1 0 189000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_46
timestamp 1765222618
transform 1 0 213000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_47
timestamp 1765222618
transform 1 0 211000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_48
timestamp 1765222618
transform 1 0 209000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_49
timestamp 1765222618
transform 1 0 207000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_50
timestamp 1765222618
transform 1 0 205000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_51
timestamp 1765222618
transform 1 0 203000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_52
timestamp 1765222618
transform 1 0 201000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_53
timestamp 1765222618
transform 1 0 199000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_54
timestamp 1765222618
transform 1 0 197000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_55
timestamp 1765222618
transform 1 0 195000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_56
timestamp 1765222618
transform 1 0 193000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_57
timestamp 1765222618
transform 1 0 191000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_58
timestamp 1765222618
transform 1 0 246000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_60
timestamp 1765222618
transform 1 0 232000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_61
timestamp 1765222618
transform 1 0 234000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_62
timestamp 1765222618
transform 1 0 236000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_63
timestamp 1765222618
transform 1 0 238000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_64
timestamp 1765222618
transform 1 0 240000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_65
timestamp 1765222618
transform 1 0 242000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_66
timestamp 1765222618
transform 1 0 244000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_67
timestamp 1765222618
transform 1 0 268000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_68
timestamp 1765222618
transform 1 0 266000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_69
timestamp 1765222618
transform 1 0 264000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_70
timestamp 1765222618
transform 1 0 262000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_71
timestamp 1765222618
transform 1 0 260000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_72
timestamp 1765222618
transform 1 0 258000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_73
timestamp 1765222618
transform 1 0 256000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_74
timestamp 1765222618
transform 1 0 254000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_75
timestamp 1765222618
transform 1 0 252000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_76
timestamp 1765222618
transform 1 0 250000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_77
timestamp 1765222618
transform 1 0 248000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_78
timestamp 1765222618
transform 1 0 303000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_79
timestamp 1765222618
transform 1 0 301000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_80
timestamp 1765222618
transform 1 0 285000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_81
timestamp 1765222618
transform 1 0 287000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_82
timestamp 1765222618
transform 1 0 289000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_83
timestamp 1765222618
transform 1 0 291000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_84
timestamp 1765222618
transform 1 0 293000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_85
timestamp 1765222618
transform 1 0 295000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_86
timestamp 1765222618
transform 1 0 297000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_87
timestamp 1765222618
transform 1 0 299000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_88
timestamp 1765222618
transform 1 0 323000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_89
timestamp 1765222618
transform 1 0 321000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_90
timestamp 1765222618
transform 1 0 319000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_91
timestamp 1765222618
transform 1 0 317000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_92
timestamp 1765222618
transform 1 0 315000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_93
timestamp 1765222618
transform 1 0 313000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_94
timestamp 1765222618
transform 1 0 311000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_95
timestamp 1765222618
transform 1 0 309000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_96
timestamp 1765222618
transform 1 0 307000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_97
timestamp 1765222618
transform 1 0 305000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_98
timestamp 1765222618
transform 1 0 360000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_99
timestamp 1765222618
transform 1 0 358000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_100
timestamp 1765222618
transform 1 0 356000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_102
timestamp 1765222618
transform 1 0 342000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_103
timestamp 1765222618
transform 1 0 344000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_104
timestamp 1765222618
transform 1 0 346000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_105
timestamp 1765222618
transform 1 0 348000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_106
timestamp 1765222618
transform 1 0 350000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_107
timestamp 1765222618
transform 1 0 352000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_108
timestamp 1765222618
transform 1 0 354000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_109
timestamp 1765222618
transform 1 0 378000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_110
timestamp 1765222618
transform 1 0 376000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_111
timestamp 1765222618
transform 1 0 374000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_112
timestamp 1765222618
transform 1 0 372000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_113
timestamp 1765222618
transform 1 0 370000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_114
timestamp 1765222618
transform 1 0 368000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_115
timestamp 1765222618
transform 1 0 366000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_116
timestamp 1765222618
transform 1 0 364000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_117
timestamp 1765222618
transform 1 0 362000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_118
timestamp 1765222618
transform 1 0 415000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_119
timestamp 1765222618
transform 1 0 413000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_120
timestamp 1765222618
transform 1 0 411000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_122
timestamp 1765222618
transform 1 0 397000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_123
timestamp 1765222618
transform 1 0 399000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_124
timestamp 1765222618
transform 1 0 401000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_125
timestamp 1765222618
transform 1 0 403000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_126
timestamp 1765222618
transform 1 0 405000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_127
timestamp 1765222618
transform 1 0 407000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_128
timestamp 1765222618
transform 1 0 409000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_129
timestamp 1765222618
transform 1 0 433000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_130
timestamp 1765222618
transform 1 0 431000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_131
timestamp 1765222618
transform 1 0 429000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_132
timestamp 1765222618
transform 1 0 427000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_133
timestamp 1765222618
transform 1 0 425000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_134
timestamp 1765222618
transform 1 0 423000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_135
timestamp 1765222618
transform 1 0 421000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_136
timestamp 1765222618
transform 1 0 419000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_137
timestamp 1765222618
transform 1 0 417000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_139
timestamp 1765222618
transform 1 0 452000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_140
timestamp 1765222618
transform 1 0 454000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_141
timestamp 1765222618
transform 1 0 456000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_142
timestamp 1765222618
transform 1 0 458000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_143
timestamp 1765222618
transform 1 0 460000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_144
timestamp 1765222618
transform 1 0 462000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_145
timestamp 1765222618
transform 1 0 466000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_146
timestamp 1765222618
transform 1 0 464000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_147
timestamp 1765222618
transform 1 0 470000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_148
timestamp 1765222618
transform 1 0 468000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_149
timestamp 1765222618
transform 1 0 474000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_150
timestamp 1765222618
transform 1 0 472000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_151
timestamp 1765222618
transform 1 0 478000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_152
timestamp 1765222618
transform 1 0 476000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_153
timestamp 1765222618
transform 1 0 482000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_154
timestamp 1765222618
transform 1 0 480000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_155
timestamp 1765222618
transform 1 0 486000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_156
timestamp 1765222618
transform 1 0 484000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_157
timestamp 1765222618
transform 1 0 488000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_175
timestamp 1765222618
transform 1 0 541000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_176
timestamp 1765222618
transform 1 0 539000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_177
timestamp 1765222618
transform 1 0 543000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_179
timestamp 1765222618
transform 1 0 562000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_180
timestamp 1765222618
transform 1 0 564000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_181
timestamp 1765222618
transform 1 0 566000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_182
timestamp 1765222618
transform 1 0 568000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_183
timestamp 1765222618
transform 1 0 570000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_184
timestamp 1765222618
transform 1 0 572000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_185
timestamp 1765222618
transform 1 0 576000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_186
timestamp 1765222618
transform 1 0 574000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_187
timestamp 1765222618
transform 1 0 580000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_188
timestamp 1765222618
transform 1 0 578000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_189
timestamp 1765222618
transform 1 0 584000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_190
timestamp 1765222618
transform 1 0 582000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_191
timestamp 1765222618
transform 1 0 588000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_192
timestamp 1765222618
transform 1 0 586000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_195
timestamp 1765222618
transform 1 0 596000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_196
timestamp 1765222618
transform 1 0 594000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_197
timestamp 1765222618
transform 1 0 598000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_198
timestamp 1765222618
transform 1 0 615000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_199
timestamp 1765222618
transform 1 0 617000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_200
timestamp 1765222618
transform 1 0 619000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_201
timestamp 1765222618
transform 1 0 621000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_202
timestamp 1765222618
transform 1 0 623000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_203
timestamp 1765222618
transform 1 0 625000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_204
timestamp 1765222618
transform 1 0 627000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_205
timestamp 1765222618
transform 1 0 631000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_206
timestamp 1765222618
transform 1 0 629000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_207
timestamp 1765222618
transform 1 0 635000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_208
timestamp 1765222618
transform 1 0 633000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_209
timestamp 1765222618
transform 1 0 639000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_210
timestamp 1765222618
transform 1 0 637000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_211
timestamp 1765222618
transform 1 0 643000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_212
timestamp 1765222618
transform 1 0 641000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_213
timestamp 1765222618
transform 1 0 647000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_214
timestamp 1765222618
transform 1 0 645000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_215
timestamp 1765222618
transform 1 0 651000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_216
timestamp 1765222618
transform 1 0 649000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_217
timestamp 1765222618
transform 1 0 653000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_218
timestamp 1765222618
transform 1 0 670000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_219
timestamp 1765222618
transform 1 0 672000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_220
timestamp 1765222618
transform 1 0 674000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_221
timestamp 1765222618
transform 1 0 676000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_222
timestamp 1765222618
transform 1 0 678000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_223
timestamp 1765222618
transform 1 0 680000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_224
timestamp 1765222618
transform 1 0 682000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_225
timestamp 1765222618
transform 1 0 686000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_226
timestamp 1765222618
transform 1 0 684000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_227
timestamp 1765222618
transform 1 0 690000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_228
timestamp 1765222618
transform 1 0 688000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_229
timestamp 1765222618
transform 1 0 694000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_230
timestamp 1765222618
transform 1 0 692000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_231
timestamp 1765222618
transform 1 0 698000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_232
timestamp 1765222618
transform 1 0 696000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_233
timestamp 1765222618
transform 1 0 702000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_234
timestamp 1765222618
transform 1 0 700000 0 1 0
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_238
timestamp 1765222618
transform 0 -1 776000 1 0 71000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_239
timestamp 1765222618
transform 0 -1 776000 1 0 73000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_240
timestamp 1765222618
transform 0 -1 776000 1 0 75000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_241
timestamp 1765222618
transform 0 -1 776000 1 0 77000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_242
timestamp 1765222618
transform 0 -1 776000 1 0 79000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_243
timestamp 1765222618
transform 0 -1 776000 1 0 81000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_244
timestamp 1765222618
transform 0 -1 776000 1 0 83000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_245
timestamp 1765222618
transform 0 -1 776000 1 0 85000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_246
timestamp 1765222618
transform 0 -1 776000 1 0 87000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_247
timestamp 1765222618
transform 0 -1 776000 1 0 112000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_248
timestamp 1765222618
transform 0 -1 776000 1 0 108000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_249
timestamp 1765222618
transform 0 -1 776000 1 0 110000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_250
timestamp 1765222618
transform 0 -1 776000 1 0 116000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_251
timestamp 1765222618
transform 0 -1 776000 1 0 114000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_252
timestamp 1765222618
transform 0 -1 776000 1 0 120000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_253
timestamp 1765222618
transform 0 -1 776000 1 0 118000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_254
timestamp 1765222618
transform 0 -1 776000 1 0 124000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_255
timestamp 1765222618
transform 0 -1 776000 1 0 122000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_256
timestamp 1765222618
transform 0 -1 776000 1 0 128000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_257
timestamp 1765222618
transform 0 -1 776000 1 0 126000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_258
timestamp 1765222618
transform 0 -1 776000 1 0 130000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_259
timestamp 1765222618
transform 0 -1 776000 1 0 106000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_262
timestamp 1765222618
transform 0 -1 776000 1 0 149000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_263
timestamp 1765222618
transform 0 -1 776000 1 0 151000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_264
timestamp 1765222618
transform 0 -1 776000 1 0 153000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_265
timestamp 1765222618
transform 0 -1 776000 1 0 157000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_266
timestamp 1765222618
transform 0 -1 776000 1 0 155000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_267
timestamp 1765222618
transform 0 -1 776000 1 0 161000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_268
timestamp 1765222618
transform 0 -1 776000 1 0 159000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_269
timestamp 1765222618
transform 0 -1 776000 1 0 165000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_270
timestamp 1765222618
transform 0 -1 776000 1 0 163000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_271
timestamp 1765222618
transform 0 -1 776000 1 0 169000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_272
timestamp 1765222618
transform 0 -1 776000 1 0 167000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_273
timestamp 1765222618
transform 0 -1 776000 1 0 173000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_274
timestamp 1765222618
transform 0 -1 776000 1 0 171000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_276
timestamp 1765222618
transform 0 -1 776000 1 0 192000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_277
timestamp 1765222618
transform 0 -1 776000 1 0 194000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_278
timestamp 1765222618
transform 0 -1 776000 1 0 196000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_279
timestamp 1765222618
transform 0 -1 776000 1 0 200000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_280
timestamp 1765222618
transform 0 -1 776000 1 0 198000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_281
timestamp 1765222618
transform 0 -1 776000 1 0 204000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_282
timestamp 1765222618
transform 0 -1 776000 1 0 202000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_283
timestamp 1765222618
transform 0 -1 776000 1 0 208000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_284
timestamp 1765222618
transform 0 -1 776000 1 0 206000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_285
timestamp 1765222618
transform 0 -1 776000 1 0 212000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_286
timestamp 1765222618
transform 0 -1 776000 1 0 210000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_287
timestamp 1765222618
transform 0 -1 776000 1 0 216000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_288
timestamp 1765222618
transform 0 -1 776000 1 0 214000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_290
timestamp 1765222618
transform 0 -1 776000 1 0 235000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_291
timestamp 1765222618
transform 0 -1 776000 1 0 237000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_292
timestamp 1765222618
transform 0 -1 776000 1 0 239000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_293
timestamp 1765222618
transform 0 -1 776000 1 0 243000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_294
timestamp 1765222618
transform 0 -1 776000 1 0 241000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_295
timestamp 1765222618
transform 0 -1 776000 1 0 247000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_296
timestamp 1765222618
transform 0 -1 776000 1 0 245000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_297
timestamp 1765222618
transform 0 -1 776000 1 0 251000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_298
timestamp 1765222618
transform 0 -1 776000 1 0 249000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_299
timestamp 1765222618
transform 0 -1 776000 1 0 255000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_300
timestamp 1765222618
transform 0 -1 776000 1 0 253000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_301
timestamp 1765222618
transform 0 -1 776000 1 0 259000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_302
timestamp 1765222618
transform 0 -1 776000 1 0 257000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_304
timestamp 1765222618
transform 0 -1 776000 1 0 278000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_305
timestamp 1765222618
transform 0 -1 776000 1 0 280000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_306
timestamp 1765222618
transform 0 -1 776000 1 0 282000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_307
timestamp 1765222618
transform 0 -1 776000 1 0 286000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_308
timestamp 1765222618
transform 0 -1 776000 1 0 284000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_309
timestamp 1765222618
transform 0 -1 776000 1 0 290000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_310
timestamp 1765222618
transform 0 -1 776000 1 0 288000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_311
timestamp 1765222618
transform 0 -1 776000 1 0 294000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_312
timestamp 1765222618
transform 0 -1 776000 1 0 292000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_313
timestamp 1765222618
transform 0 -1 776000 1 0 298000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_314
timestamp 1765222618
transform 0 -1 776000 1 0 296000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_315
timestamp 1765222618
transform 0 -1 776000 1 0 302000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_316
timestamp 1765222618
transform 0 -1 776000 1 0 300000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_318
timestamp 1765222618
transform 0 -1 776000 1 0 321000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_319
timestamp 1765222618
transform 0 -1 776000 1 0 323000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_320
timestamp 1765222618
transform 0 -1 776000 1 0 325000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_321
timestamp 1765222618
transform 0 -1 776000 1 0 329000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_322
timestamp 1765222618
transform 0 -1 776000 1 0 327000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_323
timestamp 1765222618
transform 0 -1 776000 1 0 333000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_324
timestamp 1765222618
transform 0 -1 776000 1 0 331000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_325
timestamp 1765222618
transform 0 -1 776000 1 0 337000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_326
timestamp 1765222618
transform 0 -1 776000 1 0 335000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_327
timestamp 1765222618
transform 0 -1 776000 1 0 341000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_328
timestamp 1765222618
transform 0 -1 776000 1 0 339000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_329
timestamp 1765222618
transform 0 -1 776000 1 0 345000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_330
timestamp 1765222618
transform 0 -1 776000 1 0 343000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_332
timestamp 1765222618
transform 0 -1 776000 1 0 364000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_333
timestamp 1765222618
transform 0 -1 776000 1 0 366000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_334
timestamp 1765222618
transform 0 -1 776000 1 0 368000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_335
timestamp 1765222618
transform 0 -1 776000 1 0 372000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_336
timestamp 1765222618
transform 0 -1 776000 1 0 370000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_337
timestamp 1765222618
transform 0 -1 776000 1 0 376000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_338
timestamp 1765222618
transform 0 -1 776000 1 0 374000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_339
timestamp 1765222618
transform 0 -1 776000 1 0 380000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_340
timestamp 1765222618
transform 0 -1 776000 1 0 378000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_341
timestamp 1765222618
transform 0 -1 776000 1 0 384000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_342
timestamp 1765222618
transform 0 -1 776000 1 0 382000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_343
timestamp 1765222618
transform 0 -1 776000 1 0 388000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_344
timestamp 1765222618
transform 0 -1 776000 1 0 386000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_345
timestamp 1765222618
transform 0 -1 776000 1 0 405000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_346
timestamp 1765222618
transform 0 -1 776000 1 0 407000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_347
timestamp 1765222618
transform 0 -1 776000 1 0 409000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_348
timestamp 1765222618
transform 0 -1 776000 1 0 411000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_349
timestamp 1765222618
transform 0 -1 776000 1 0 415000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_350
timestamp 1765222618
transform 0 -1 776000 1 0 413000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_351
timestamp 1765222618
transform 0 -1 776000 1 0 419000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_352
timestamp 1765222618
transform 0 -1 776000 1 0 417000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_353
timestamp 1765222618
transform 0 -1 776000 1 0 423000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_354
timestamp 1765222618
transform 0 -1 776000 1 0 421000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_355
timestamp 1765222618
transform 0 -1 776000 1 0 427000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_356
timestamp 1765222618
transform 0 -1 776000 1 0 425000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_357
timestamp 1765222618
transform 0 -1 776000 1 0 431000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_358
timestamp 1765222618
transform 0 -1 776000 1 0 429000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_359
timestamp 1765222618
transform 0 -1 776000 1 0 448000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_360
timestamp 1765222618
transform 0 -1 776000 1 0 450000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_361
timestamp 1765222618
transform 0 -1 776000 1 0 452000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_362
timestamp 1765222618
transform 0 -1 776000 1 0 454000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_363
timestamp 1765222618
transform 0 -1 776000 1 0 458000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_364
timestamp 1765222618
transform 0 -1 776000 1 0 456000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_365
timestamp 1765222618
transform 0 -1 776000 1 0 462000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_366
timestamp 1765222618
transform 0 -1 776000 1 0 460000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_367
timestamp 1765222618
transform 0 -1 776000 1 0 466000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_368
timestamp 1765222618
transform 0 -1 776000 1 0 464000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_369
timestamp 1765222618
transform 0 -1 776000 1 0 470000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_370
timestamp 1765222618
transform 0 -1 776000 1 0 468000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_371
timestamp 1765222618
transform 0 -1 776000 1 0 474000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_372
timestamp 1765222618
transform 0 -1 776000 1 0 472000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_373
timestamp 1765222618
transform 0 -1 776000 1 0 491000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_374
timestamp 1765222618
transform 0 -1 776000 1 0 493000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_375
timestamp 1765222618
transform 0 -1 776000 1 0 495000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_376
timestamp 1765222618
transform 0 -1 776000 1 0 497000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_377
timestamp 1765222618
transform 0 -1 776000 1 0 501000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_378
timestamp 1765222618
transform 0 -1 776000 1 0 499000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_379
timestamp 1765222618
transform 0 -1 776000 1 0 505000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_380
timestamp 1765222618
transform 0 -1 776000 1 0 503000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_381
timestamp 1765222618
transform 0 -1 776000 1 0 509000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_382
timestamp 1765222618
transform 0 -1 776000 1 0 507000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_383
timestamp 1765222618
transform 0 -1 776000 1 0 513000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_384
timestamp 1765222618
transform 0 -1 776000 1 0 511000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_385
timestamp 1765222618
transform 0 -1 776000 1 0 517000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_386
timestamp 1765222618
transform 0 -1 776000 1 0 515000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_388
timestamp 1765222618
transform 0 -1 776000 1 0 536000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_389
timestamp 1765222618
transform 0 -1 776000 1 0 538000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_390
timestamp 1765222618
transform 0 -1 776000 1 0 540000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_391
timestamp 1765222618
transform 0 -1 776000 1 0 544000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_392
timestamp 1765222618
transform 0 -1 776000 1 0 542000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_393
timestamp 1765222618
transform 0 -1 776000 1 0 548000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_394
timestamp 1765222618
transform 0 -1 776000 1 0 546000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_395
timestamp 1765222618
transform 0 -1 776000 1 0 552000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_396
timestamp 1765222618
transform 0 -1 776000 1 0 550000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_397
timestamp 1765222618
transform 0 -1 776000 1 0 556000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_398
timestamp 1765222618
transform 0 -1 776000 1 0 554000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_399
timestamp 1765222618
transform 0 -1 776000 1 0 560000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_400
timestamp 1765222618
transform 0 -1 776000 1 0 558000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_402
timestamp 1765222618
transform 0 -1 776000 1 0 579000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_403
timestamp 1765222618
transform 0 -1 776000 1 0 581000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_404
timestamp 1765222618
transform 0 -1 776000 1 0 583000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_405
timestamp 1765222618
transform 0 -1 776000 1 0 587000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_406
timestamp 1765222618
transform 0 -1 776000 1 0 585000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_407
timestamp 1765222618
transform 0 -1 776000 1 0 591000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_408
timestamp 1765222618
transform 0 -1 776000 1 0 589000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_409
timestamp 1765222618
transform 0 -1 776000 1 0 595000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_410
timestamp 1765222618
transform 0 -1 776000 1 0 593000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_411
timestamp 1765222618
transform 0 -1 776000 1 0 599000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_412
timestamp 1765222618
transform 0 -1 776000 1 0 597000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_413
timestamp 1765222618
transform 0 -1 776000 1 0 603000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_414
timestamp 1765222618
transform 0 -1 776000 1 0 601000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_416
timestamp 1765222618
transform 0 -1 776000 1 0 622000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_417
timestamp 1765222618
transform 0 -1 776000 1 0 624000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_418
timestamp 1765222618
transform 0 -1 776000 1 0 626000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_419
timestamp 1765222618
transform 0 -1 776000 1 0 630000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_420
timestamp 1765222618
transform 0 -1 776000 1 0 628000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_421
timestamp 1765222618
transform 0 -1 776000 1 0 634000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_422
timestamp 1765222618
transform 0 -1 776000 1 0 632000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_423
timestamp 1765222618
transform 0 -1 776000 1 0 638000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_424
timestamp 1765222618
transform 0 -1 776000 1 0 636000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_425
timestamp 1765222618
transform 0 -1 776000 1 0 642000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_426
timestamp 1765222618
transform 0 -1 776000 1 0 640000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_427
timestamp 1765222618
transform 0 -1 776000 1 0 646000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_428
timestamp 1765222618
transform 0 -1 776000 1 0 644000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_430
timestamp 1765222618
transform 0 -1 776000 1 0 665000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_431
timestamp 1765222618
transform 0 -1 776000 1 0 667000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_432
timestamp 1765222618
transform 0 -1 776000 1 0 669000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_433
timestamp 1765222618
transform 0 -1 776000 1 0 673000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_434
timestamp 1765222618
transform 0 -1 776000 1 0 671000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_435
timestamp 1765222618
transform 0 -1 776000 1 0 677000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_436
timestamp 1765222618
transform 0 -1 776000 1 0 675000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_437
timestamp 1765222618
transform 0 -1 776000 1 0 681000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_438
timestamp 1765222618
transform 0 -1 776000 1 0 679000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_439
timestamp 1765222618
transform 0 -1 776000 1 0 685000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_440
timestamp 1765222618
transform 0 -1 776000 1 0 683000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_441
timestamp 1765222618
transform 0 -1 776000 1 0 689000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_442
timestamp 1765222618
transform 0 -1 776000 1 0 687000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_444
timestamp 1765222618
transform 0 -1 776000 1 0 708000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_445
timestamp 1765222618
transform 0 -1 776000 1 0 710000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_446
timestamp 1765222618
transform 0 -1 776000 1 0 712000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_447
timestamp 1765222618
transform 0 -1 776000 1 0 716000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_448
timestamp 1765222618
transform 0 -1 776000 1 0 714000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_449
timestamp 1765222618
transform 0 -1 776000 1 0 720000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_450
timestamp 1765222618
transform 0 -1 776000 1 0 718000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_451
timestamp 1765222618
transform 0 -1 776000 1 0 724000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_452
timestamp 1765222618
transform 0 -1 776000 1 0 722000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_453
timestamp 1765222618
transform 0 -1 776000 1 0 728000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_454
timestamp 1765222618
transform 0 -1 776000 1 0 726000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_455
timestamp 1765222618
transform 0 -1 776000 1 0 732000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_456
timestamp 1765222618
transform 0 -1 776000 1 0 730000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_458
timestamp 1765222618
transform 0 -1 776000 1 0 751000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_459
timestamp 1765222618
transform 0 -1 776000 1 0 753000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_460
timestamp 1765222618
transform 0 -1 776000 1 0 755000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_461
timestamp 1765222618
transform 0 -1 776000 1 0 759000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_462
timestamp 1765222618
transform 0 -1 776000 1 0 757000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_463
timestamp 1765222618
transform 0 -1 776000 1 0 763000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_464
timestamp 1765222618
transform 0 -1 776000 1 0 761000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_465
timestamp 1765222618
transform 0 -1 776000 1 0 767000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_466
timestamp 1765222618
transform 0 -1 776000 1 0 765000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_467
timestamp 1765222618
transform 0 -1 776000 1 0 771000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_468
timestamp 1765222618
transform 0 -1 776000 1 0 769000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_469
timestamp 1765222618
transform 0 -1 776000 1 0 775000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_470
timestamp 1765222618
transform 0 -1 776000 1 0 773000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_471
timestamp 1765222618
transform 0 -1 776000 1 0 792000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_472
timestamp 1765222618
transform 0 -1 776000 1 0 794000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_473
timestamp 1765222618
transform 0 -1 776000 1 0 796000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_474
timestamp 1765222618
transform 0 -1 776000 1 0 798000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_475
timestamp 1765222618
transform 0 -1 776000 1 0 802000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_476
timestamp 1765222618
transform 0 -1 776000 1 0 800000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_477
timestamp 1765222618
transform 0 -1 776000 1 0 806000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_478
timestamp 1765222618
transform 0 -1 776000 1 0 804000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_479
timestamp 1765222618
transform 0 -1 776000 1 0 810000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_480
timestamp 1765222618
transform 0 -1 776000 1 0 808000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_481
timestamp 1765222618
transform 0 -1 776000 1 0 814000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_482
timestamp 1765222618
transform 0 -1 776000 1 0 812000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_483
timestamp 1765222618
transform 0 -1 776000 1 0 818000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_484
timestamp 1765222618
transform 0 -1 776000 1 0 816000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_486
timestamp 1765222618
transform 0 -1 776000 1 0 837000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_487
timestamp 1765222618
transform 0 -1 776000 1 0 839000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_488
timestamp 1765222618
transform 0 -1 776000 1 0 841000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_489
timestamp 1765222618
transform 0 -1 776000 1 0 845000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_490
timestamp 1765222618
transform 0 -1 776000 1 0 843000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_491
timestamp 1765222618
transform 0 -1 776000 1 0 849000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_492
timestamp 1765222618
transform 0 -1 776000 1 0 847000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_493
timestamp 1765222618
transform 0 -1 776000 1 0 853000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_494
timestamp 1765222618
transform 0 -1 776000 1 0 851000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_495
timestamp 1765222618
transform 0 -1 776000 1 0 857000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_496
timestamp 1765222618
transform 0 -1 776000 1 0 855000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_497
timestamp 1765222618
transform 0 -1 776000 1 0 861000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_498
timestamp 1765222618
transform 0 -1 776000 1 0 859000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_499
timestamp 1765222618
transform 0 -1 776000 1 0 878000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_500
timestamp 1765222618
transform 0 -1 776000 1 0 880000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_501
timestamp 1765222618
transform 0 -1 776000 1 0 882000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_502
timestamp 1765222618
transform 0 -1 776000 1 0 884000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_503
timestamp 1765222618
transform 0 -1 776000 1 0 888000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_504
timestamp 1765222618
transform 0 -1 776000 1 0 886000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_505
timestamp 1765222618
transform 0 -1 776000 1 0 892000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_506
timestamp 1765222618
transform 0 -1 776000 1 0 890000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_507
timestamp 1765222618
transform 0 -1 776000 1 0 896000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_508
timestamp 1765222618
transform 0 -1 776000 1 0 894000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_509
timestamp 1765222618
transform 0 -1 776000 1 0 900000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_510
timestamp 1765222618
transform 0 -1 776000 1 0 898000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_511
timestamp 1765222618
transform 0 -1 776000 1 0 904000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_512
timestamp 1765222618
transform 0 -1 776000 1 0 902000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_513
timestamp 1765222618
transform 0 -1 776000 1 0 925000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_515
timestamp 1765222618
transform 0 -1 776000 1 0 923000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_516
timestamp 1765222618
transform 0 -1 776000 1 0 929000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_517
timestamp 1765222618
transform 0 -1 776000 1 0 927000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_518
timestamp 1765222618
transform 0 -1 776000 1 0 933000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_519
timestamp 1765222618
transform 0 -1 776000 1 0 931000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_520
timestamp 1765222618
transform 0 -1 776000 1 0 937000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_521
timestamp 1765222618
transform 0 -1 776000 1 0 935000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_522
timestamp 1765222618
transform 0 -1 776000 1 0 941000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_523
timestamp 1765222618
transform 0 -1 776000 1 0 939000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_524
timestamp 1765222618
transform -1 0 693000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_525
timestamp 1765222618
transform -1 0 695000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_526
timestamp 1765222618
transform -1 0 705000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_527
timestamp 1765222618
transform -1 0 703000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_528
timestamp 1765222618
transform -1 0 701000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_529
timestamp 1765222618
transform -1 0 699000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_530
timestamp 1765222618
transform -1 0 697000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_531
timestamp 1765222618
transform -1 0 677000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_532
timestamp 1765222618
transform -1 0 679000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_533
timestamp 1765222618
transform -1 0 681000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_534
timestamp 1765222618
transform -1 0 683000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_535
timestamp 1765222618
transform -1 0 685000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_536
timestamp 1765222618
transform -1 0 687000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_537
timestamp 1765222618
transform -1 0 691000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_538
timestamp 1765222618
transform -1 0 689000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_539
timestamp 1765222618
transform -1 0 675000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_540
timestamp 1765222618
transform -1 0 673000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_541
timestamp 1765222618
transform -1 0 671000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_542
timestamp 1765222618
transform -1 0 652000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_543
timestamp 1765222618
transform -1 0 650000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_544
timestamp 1765222618
transform -1 0 648000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_546
timestamp 1765222618
transform -1 0 636000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_547
timestamp 1765222618
transform -1 0 634000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_548
timestamp 1765222618
transform -1 0 632000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_549
timestamp 1765222618
transform -1 0 644000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_550
timestamp 1765222618
transform -1 0 642000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_551
timestamp 1765222618
transform -1 0 640000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_552
timestamp 1765222618
transform -1 0 638000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_553
timestamp 1765222618
transform -1 0 646000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_554
timestamp 1765222618
transform -1 0 622000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_555
timestamp 1765222618
transform -1 0 620000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_556
timestamp 1765222618
transform -1 0 618000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_557
timestamp 1765222618
transform -1 0 630000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_558
timestamp 1765222618
transform -1 0 628000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_559
timestamp 1765222618
transform -1 0 626000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_560
timestamp 1765222618
transform -1 0 624000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_561
timestamp 1765222618
transform -1 0 616000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_562
timestamp 1765222618
transform -1 0 587000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_563
timestamp 1765222618
transform -1 0 589000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_564
timestamp 1765222618
transform -1 0 591000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_565
timestamp 1765222618
transform -1 0 593000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_566
timestamp 1765222618
transform -1 0 595000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_567
timestamp 1765222618
transform -1 0 597000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_568
timestamp 1765222618
transform -1 0 599000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_569
timestamp 1765222618
transform -1 0 575000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_570
timestamp 1765222618
transform -1 0 573000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_571
timestamp 1765222618
transform -1 0 581000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_572
timestamp 1765222618
transform -1 0 579000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_573
timestamp 1765222618
transform -1 0 577000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_574
timestamp 1765222618
transform -1 0 583000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_575
timestamp 1765222618
transform -1 0 585000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_576
timestamp 1765222618
transform -1 0 565000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_577
timestamp 1765222618
transform -1 0 563000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_578
timestamp 1765222618
transform -1 0 561000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_579
timestamp 1765222618
transform -1 0 571000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_580
timestamp 1765222618
transform -1 0 569000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_581
timestamp 1765222618
transform -1 0 567000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_583
timestamp 1765222618
transform -1 0 542000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_584
timestamp 1765222618
transform -1 0 528000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_585
timestamp 1765222618
transform -1 0 530000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_586
timestamp 1765222618
transform -1 0 526000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_587
timestamp 1765222618
transform -1 0 536000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_588
timestamp 1765222618
transform -1 0 534000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_589
timestamp 1765222618
transform -1 0 532000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_590
timestamp 1765222618
transform -1 0 540000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_591
timestamp 1765222618
transform -1 0 538000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_592
timestamp 1765222618
transform -1 0 512000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_593
timestamp 1765222618
transform -1 0 514000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_594
timestamp 1765222618
transform -1 0 516000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_595
timestamp 1765222618
transform -1 0 518000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_596
timestamp 1765222618
transform -1 0 520000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_597
timestamp 1765222618
transform -1 0 522000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_598
timestamp 1765222618
transform -1 0 524000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_599
timestamp 1765222618
transform -1 0 506000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_600
timestamp 1765222618
transform -1 0 508000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_601
timestamp 1765222618
transform -1 0 510000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_602
timestamp 1765222618
transform -1 0 483000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_603
timestamp 1765222618
transform -1 0 481000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_604
timestamp 1765222618
transform -1 0 485000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_605
timestamp 1765222618
transform -1 0 487000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_607
timestamp 1765222618
transform -1 0 467000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_608
timestamp 1765222618
transform -1 0 469000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_609
timestamp 1765222618
transform -1 0 471000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_610
timestamp 1765222618
transform -1 0 473000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_611
timestamp 1765222618
transform -1 0 475000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_612
timestamp 1765222618
transform -1 0 477000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_613
timestamp 1765222618
transform -1 0 479000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_614
timestamp 1765222618
transform -1 0 453000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_615
timestamp 1765222618
transform -1 0 451000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_616
timestamp 1765222618
transform -1 0 461000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_617
timestamp 1765222618
transform -1 0 459000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_618
timestamp 1765222618
transform -1 0 457000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_619
timestamp 1765222618
transform -1 0 455000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_620
timestamp 1765222618
transform -1 0 463000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_621
timestamp 1765222618
transform -1 0 465000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_622
timestamp 1765222618
transform -1 0 422000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_623
timestamp 1765222618
transform -1 0 424000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_624
timestamp 1765222618
transform -1 0 426000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_625
timestamp 1765222618
transform -1 0 428000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_626
timestamp 1765222618
transform -1 0 430000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_627
timestamp 1765222618
transform -1 0 432000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_629
timestamp 1765222618
transform -1 0 406000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_630
timestamp 1765222618
transform -1 0 408000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_631
timestamp 1765222618
transform -1 0 410000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_632
timestamp 1765222618
transform -1 0 412000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_633
timestamp 1765222618
transform -1 0 414000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_634
timestamp 1765222618
transform -1 0 416000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_635
timestamp 1765222618
transform -1 0 418000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_636
timestamp 1765222618
transform -1 0 420000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_637
timestamp 1765222618
transform -1 0 400000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_638
timestamp 1765222618
transform -1 0 398000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_639
timestamp 1765222618
transform -1 0 396000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_640
timestamp 1765222618
transform -1 0 402000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_641
timestamp 1765222618
transform -1 0 404000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_642
timestamp 1765222618
transform -1 0 379000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_643
timestamp 1765222618
transform -1 0 377000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_644
timestamp 1765222618
transform -1 0 365000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_645
timestamp 1765222618
transform -1 0 367000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_646
timestamp 1765222618
transform -1 0 363000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_647
timestamp 1765222618
transform -1 0 361000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_648
timestamp 1765222618
transform -1 0 369000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_649
timestamp 1765222618
transform -1 0 375000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_650
timestamp 1765222618
transform -1 0 373000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_651
timestamp 1765222618
transform -1 0 371000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_652
timestamp 1765222618
transform -1 0 353000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_653
timestamp 1765222618
transform -1 0 351000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_654
timestamp 1765222618
transform -1 0 349000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_655
timestamp 1765222618
transform -1 0 347000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_656
timestamp 1765222618
transform -1 0 357000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_657
timestamp 1765222618
transform -1 0 355000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_658
timestamp 1765222618
transform -1 0 359000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_659
timestamp 1765222618
transform -1 0 345000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_660
timestamp 1765222618
transform -1 0 343000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_661
timestamp 1765222618
transform -1 0 341000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_662
timestamp 1765222618
transform -1 0 322000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_663
timestamp 1765222618
transform -1 0 320000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_664
timestamp 1765222618
transform -1 0 318000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_665
timestamp 1765222618
transform -1 0 316000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_667
timestamp 1765222618
transform -1 0 302000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_668
timestamp 1765222618
transform -1 0 300000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_669
timestamp 1765222618
transform -1 0 306000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_670
timestamp 1765222618
transform -1 0 304000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_671
timestamp 1765222618
transform -1 0 312000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_672
timestamp 1765222618
transform -1 0 308000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_673
timestamp 1765222618
transform -1 0 310000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_674
timestamp 1765222618
transform -1 0 314000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_675
timestamp 1765222618
transform -1 0 286000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_676
timestamp 1765222618
transform -1 0 290000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_677
timestamp 1765222618
transform -1 0 288000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_678
timestamp 1765222618
transform -1 0 294000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_679
timestamp 1765222618
transform -1 0 292000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_680
timestamp 1765222618
transform -1 0 296000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_681
timestamp 1765222618
transform -1 0 298000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_682
timestamp 1765222618
transform -1 0 255000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_683
timestamp 1765222618
transform -1 0 257000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_684
timestamp 1765222618
transform -1 0 259000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_685
timestamp 1765222618
transform -1 0 261000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_686
timestamp 1765222618
transform -1 0 263000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_687
timestamp 1765222618
transform -1 0 265000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_688
timestamp 1765222618
transform -1 0 267000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_690
timestamp 1765222618
transform -1 0 241000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_691
timestamp 1765222618
transform -1 0 243000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_692
timestamp 1765222618
transform -1 0 245000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_693
timestamp 1765222618
transform -1 0 247000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_694
timestamp 1765222618
transform -1 0 251000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_695
timestamp 1765222618
transform -1 0 249000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_696
timestamp 1765222618
transform -1 0 253000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_697
timestamp 1765222618
transform -1 0 237000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_698
timestamp 1765222618
transform -1 0 239000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_699
timestamp 1765222618
transform -1 0 233000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_700
timestamp 1765222618
transform -1 0 235000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_701
timestamp 1765222618
transform -1 0 231000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_702
timestamp 1765222618
transform -1 0 210000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_703
timestamp 1765222618
transform -1 0 212000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_705
timestamp 1765222618
transform -1 0 196000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_706
timestamp 1765222618
transform -1 0 208000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_707
timestamp 1765222618
transform -1 0 206000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_708
timestamp 1765222618
transform -1 0 204000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_709
timestamp 1765222618
transform -1 0 202000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_710
timestamp 1765222618
transform -1 0 198000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_711
timestamp 1765222618
transform -1 0 200000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_712
timestamp 1765222618
transform -1 0 180000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_713
timestamp 1765222618
transform -1 0 182000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_714
timestamp 1765222618
transform -1 0 194000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_715
timestamp 1765222618
transform -1 0 190000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_716
timestamp 1765222618
transform -1 0 192000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_717
timestamp 1765222618
transform -1 0 186000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_718
timestamp 1765222618
transform -1 0 188000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_719
timestamp 1765222618
transform -1 0 184000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_720
timestamp 1765222618
transform -1 0 178000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_721
timestamp 1765222618
transform -1 0 176000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_722
timestamp 1765222618
transform -1 0 151000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_723
timestamp 1765222618
transform -1 0 155000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_724
timestamp 1765222618
transform -1 0 153000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_726
timestamp 1765222618
transform -1 0 157000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_727
timestamp 1765222618
transform -1 0 139000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_728
timestamp 1765222618
transform -1 0 135000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_729
timestamp 1765222618
transform -1 0 137000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_730
timestamp 1765222618
transform -1 0 141000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_731
timestamp 1765222618
transform -1 0 149000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_732
timestamp 1765222618
transform -1 0 147000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_733
timestamp 1765222618
transform -1 0 143000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_734
timestamp 1765222618
transform -1 0 145000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_735
timestamp 1765222618
transform -1 0 123000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_736
timestamp 1765222618
transform -1 0 125000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_737
timestamp 1765222618
transform -1 0 121000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_738
timestamp 1765222618
transform -1 0 131000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_739
timestamp 1765222618
transform -1 0 133000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_740
timestamp 1765222618
transform -1 0 127000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_741
timestamp 1765222618
transform -1 0 129000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_742
timestamp 1765222618
transform -1 0 90000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_743
timestamp 1765222618
transform -1 0 92000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_744
timestamp 1765222618
transform -1 0 94000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_745
timestamp 1765222618
transform -1 0 96000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_746
timestamp 1765222618
transform -1 0 98000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_748
timestamp 1765222618
transform -1 0 102000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_749
timestamp 1765222618
transform -1 0 100000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_750
timestamp 1765222618
transform -1 0 74000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_751
timestamp 1765222618
transform -1 0 76000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_752
timestamp 1765222618
transform -1 0 78000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_753
timestamp 1765222618
transform -1 0 80000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_754
timestamp 1765222618
transform -1 0 82000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_755
timestamp 1765222618
transform -1 0 84000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_756
timestamp 1765222618
transform -1 0 86000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_757
timestamp 1765222618
transform -1 0 88000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_759
timestamp 1765222618
transform 0 1 0 -1 0 940000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_760
timestamp 1765222618
transform 0 1 0 -1 0 942000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_761
timestamp 1765222618
transform 0 1 0 -1 0 102000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_762
timestamp 1765222618
transform 0 1 0 -1 0 934000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_763
timestamp 1765222618
transform 0 1 0 -1 0 936000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_764
timestamp 1765222618
transform 0 1 0 -1 0 938000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_765
timestamp 1765222618
transform 0 1 0 -1 0 932000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_766
timestamp 1765222618
transform 0 1 0 -1 0 928000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_767
timestamp 1765222618
transform 0 1 0 -1 0 930000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_768
timestamp 1765222618
transform 0 1 0 -1 0 922000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_769
timestamp 1765222618
transform 0 1 0 -1 0 926000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_770
timestamp 1765222618
transform 0 1 0 -1 0 924000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_771
timestamp 1765222618
transform 0 1 0 -1 0 903000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_773
timestamp 1765222618
transform 0 1 0 -1 0 104000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_774
timestamp 1765222618
transform 0 1 0 -1 0 895000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_775
timestamp 1765222618
transform 0 1 0 -1 0 893000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_776
timestamp 1765222618
transform 0 1 0 -1 0 899000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_777
timestamp 1765222618
transform 0 1 0 -1 0 901000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_778
timestamp 1765222618
transform 0 1 0 -1 0 897000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_779
timestamp 1765222618
transform 0 1 0 -1 0 889000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_780
timestamp 1765222618
transform 0 1 0 -1 0 891000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_781
timestamp 1765222618
transform 0 1 0 -1 0 881000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_782
timestamp 1765222618
transform 0 1 0 -1 0 887000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_783
timestamp 1765222618
transform 0 1 0 -1 0 883000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_784
timestamp 1765222618
transform 0 1 0 -1 0 885000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_785
timestamp 1765222618
transform 0 1 0 -1 0 106000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_786
timestamp 1765222618
transform 0 1 0 -1 0 860000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_787
timestamp 1765222618
transform 0 1 0 -1 0 862000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_788
timestamp 1765222618
transform 0 1 0 -1 0 864000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_789
timestamp 1765222618
transform 0 1 0 -1 0 854000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_790
timestamp 1765222618
transform 0 1 0 -1 0 858000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_791
timestamp 1765222618
transform 0 1 0 -1 0 856000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_792
timestamp 1765222618
transform 0 1 0 -1 0 846000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_793
timestamp 1765222618
transform 0 1 0 -1 0 850000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_794
timestamp 1765222618
transform 0 1 0 -1 0 848000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_795
timestamp 1765222618
transform 0 1 0 -1 0 852000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_796
timestamp 1765222618
transform 0 1 0 -1 0 842000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_797
timestamp 1765222618
transform 0 1 0 -1 0 840000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_798
timestamp 1765222618
transform 0 1 0 -1 0 844000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_799
timestamp 1765222618
transform 0 1 0 -1 0 817000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_800
timestamp 1765222618
transform 0 1 0 -1 0 108000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_801
timestamp 1765222618
transform 0 1 0 -1 0 823000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_802
timestamp 1765222618
transform 0 1 0 -1 0 821000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_803
timestamp 1765222618
transform 0 1 0 -1 0 819000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_804
timestamp 1765222618
transform 0 1 0 -1 0 815000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_805
timestamp 1765222618
transform 0 1 0 -1 0 811000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_806
timestamp 1765222618
transform 0 1 0 -1 0 813000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_807
timestamp 1765222618
transform 0 1 0 -1 0 809000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_808
timestamp 1765222618
transform 0 1 0 -1 0 805000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_809
timestamp 1765222618
transform 0 1 0 -1 0 803000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_810
timestamp 1765222618
transform 0 1 0 -1 0 807000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_811
timestamp 1765222618
transform 0 1 0 -1 0 801000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_812
timestamp 1765222618
transform 0 1 0 -1 0 799000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_813
timestamp 1765222618
transform 0 1 0 -1 0 776000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_814
timestamp 1765222618
transform 0 1 0 -1 0 774000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_815
timestamp 1765222618
transform 0 1 0 -1 0 778000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_816
timestamp 1765222618
transform 0 1 0 -1 0 780000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_817
timestamp 1765222618
transform 0 1 0 -1 0 782000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_818
timestamp 1765222618
transform 0 1 0 -1 0 110000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_819
timestamp 1765222618
transform 0 1 0 -1 0 772000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_820
timestamp 1765222618
transform 0 1 0 -1 0 760000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_821
timestamp 1765222618
transform 0 1 0 -1 0 764000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_822
timestamp 1765222618
transform 0 1 0 -1 0 762000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_823
timestamp 1765222618
transform 0 1 0 -1 0 768000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_824
timestamp 1765222618
transform 0 1 0 -1 0 766000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_825
timestamp 1765222618
transform 0 1 0 -1 0 770000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_826
timestamp 1765222618
transform 0 1 0 -1 0 758000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_827
timestamp 1765222618
transform 0 1 0 -1 0 112000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_829
timestamp 1765222618
transform 0 1 0 -1 0 739000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_830
timestamp 1765222618
transform 0 1 0 -1 0 737000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_831
timestamp 1765222618
transform 0 1 0 -1 0 733000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_832
timestamp 1765222618
transform 0 1 0 -1 0 735000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_833
timestamp 1765222618
transform 0 1 0 -1 0 731000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_834
timestamp 1765222618
transform 0 1 0 -1 0 729000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_835
timestamp 1765222618
transform 0 1 0 -1 0 725000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_836
timestamp 1765222618
transform 0 1 0 -1 0 727000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_837
timestamp 1765222618
transform 0 1 0 -1 0 721000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_838
timestamp 1765222618
transform 0 1 0 -1 0 723000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_839
timestamp 1765222618
transform 0 1 0 -1 0 719000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_840
timestamp 1765222618
transform 0 1 0 -1 0 717000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_842
timestamp 1765222618
transform 0 1 0 -1 0 698000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_843
timestamp 1765222618
transform 0 1 0 -1 0 696000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_844
timestamp 1765222618
transform 0 1 0 -1 0 692000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_845
timestamp 1765222618
transform 0 1 0 -1 0 694000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_846
timestamp 1765222618
transform 0 1 0 -1 0 690000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_847
timestamp 1765222618
transform 0 1 0 -1 0 114000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_848
timestamp 1765222618
transform 0 1 0 -1 0 688000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_849
timestamp 1765222618
transform 0 1 0 -1 0 684000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_850
timestamp 1765222618
transform 0 1 0 -1 0 680000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_851
timestamp 1765222618
transform 0 1 0 -1 0 682000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_852
timestamp 1765222618
transform 0 1 0 -1 0 676000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_853
timestamp 1765222618
transform 0 1 0 -1 0 678000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_854
timestamp 1765222618
transform 0 1 0 -1 0 686000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_856
timestamp 1765222618
transform 0 1 0 -1 0 116000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_857
timestamp 1765222618
transform 0 1 0 -1 0 653000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_858
timestamp 1765222618
transform 0 1 0 -1 0 651000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_859
timestamp 1765222618
transform 0 1 0 -1 0 655000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_860
timestamp 1765222618
transform 0 1 0 -1 0 657000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_861
timestamp 1765222618
transform 0 1 0 -1 0 645000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_862
timestamp 1765222618
transform 0 1 0 -1 0 649000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_863
timestamp 1765222618
transform 0 1 0 -1 0 647000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_864
timestamp 1765222618
transform 0 1 0 -1 0 637000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_865
timestamp 1765222618
transform 0 1 0 -1 0 641000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_866
timestamp 1765222618
transform 0 1 0 -1 0 639000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_867
timestamp 1765222618
transform 0 1 0 -1 0 643000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_868
timestamp 1765222618
transform 0 1 0 -1 0 635000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_869
timestamp 1765222618
transform 0 1 0 -1 0 616000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_871
timestamp 1765222618
transform 0 1 0 -1 0 118000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_872
timestamp 1765222618
transform 0 1 0 -1 0 612000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_873
timestamp 1765222618
transform 0 1 0 -1 0 610000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_874
timestamp 1765222618
transform 0 1 0 -1 0 614000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_875
timestamp 1765222618
transform 0 1 0 -1 0 608000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_876
timestamp 1765222618
transform 0 1 0 -1 0 604000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_877
timestamp 1765222618
transform 0 1 0 -1 0 602000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_878
timestamp 1765222618
transform 0 1 0 -1 0 606000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_879
timestamp 1765222618
transform 0 1 0 -1 0 596000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_880
timestamp 1765222618
transform 0 1 0 -1 0 594000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_881
timestamp 1765222618
transform 0 1 0 -1 0 600000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_882
timestamp 1765222618
transform 0 1 0 -1 0 598000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_883
timestamp 1765222618
transform 0 1 0 -1 0 573000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_884
timestamp 1765222618
transform 0 1 0 -1 0 575000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_886
timestamp 1765222618
transform 0 1 0 -1 0 120000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_887
timestamp 1765222618
transform 0 1 0 -1 0 571000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_888
timestamp 1765222618
transform 0 1 0 -1 0 569000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_889
timestamp 1765222618
transform 0 1 0 -1 0 559000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_890
timestamp 1765222618
transform 0 1 0 -1 0 563000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_891
timestamp 1765222618
transform 0 1 0 -1 0 561000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_892
timestamp 1765222618
transform 0 1 0 -1 0 565000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_893
timestamp 1765222618
transform 0 1 0 -1 0 567000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_894
timestamp 1765222618
transform 0 1 0 -1 0 555000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_895
timestamp 1765222618
transform 0 1 0 -1 0 557000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_896
timestamp 1765222618
transform 0 1 0 -1 0 553000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_897
timestamp 1765222618
transform 0 1 0 -1 0 530000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_898
timestamp 1765222618
transform 0 1 0 -1 0 532000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_899
timestamp 1765222618
transform 0 1 0 -1 0 534000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_901
timestamp 1765222618
transform 0 1 0 -1 0 122000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_902
timestamp 1765222618
transform 0 1 0 -1 0 526000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_903
timestamp 1765222618
transform 0 1 0 -1 0 528000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_904
timestamp 1765222618
transform 0 1 0 -1 0 518000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_905
timestamp 1765222618
transform 0 1 0 -1 0 516000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_906
timestamp 1765222618
transform 0 1 0 -1 0 522000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_907
timestamp 1765222618
transform 0 1 0 -1 0 520000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_908
timestamp 1765222618
transform 0 1 0 -1 0 524000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_909
timestamp 1765222618
transform 0 1 0 -1 0 512000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_910
timestamp 1765222618
transform 0 1 0 -1 0 514000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_911
timestamp 1765222618
transform 0 1 0 -1 0 489000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_912
timestamp 1765222618
transform 0 1 0 -1 0 487000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_913
timestamp 1765222618
transform 0 1 0 -1 0 491000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_914
timestamp 1765222618
transform 0 1 0 -1 0 493000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_916
timestamp 1765222618
transform 0 1 0 -1 0 124000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_917
timestamp 1765222618
transform 0 1 0 -1 0 473000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_918
timestamp 1765222618
transform 0 1 0 -1 0 477000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_919
timestamp 1765222618
transform 0 1 0 -1 0 475000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_920
timestamp 1765222618
transform 0 1 0 -1 0 481000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_921
timestamp 1765222618
transform 0 1 0 -1 0 479000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_922
timestamp 1765222618
transform 0 1 0 -1 0 483000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_923
timestamp 1765222618
transform 0 1 0 -1 0 485000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_924
timestamp 1765222618
transform 0 1 0 -1 0 471000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_925
timestamp 1765222618
transform 0 1 0 -1 0 126000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_926
timestamp 1765222618
transform 0 1 0 -1 0 454000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_927
timestamp 1765222618
transform 0 1 0 -1 0 452000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_928
timestamp 1765222618
transform 0 1 0 -1 0 450000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_929
timestamp 1765222618
transform 0 1 0 -1 0 448000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_930
timestamp 1765222618
transform 0 1 0 -1 0 444000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_931
timestamp 1765222618
transform 0 1 0 -1 0 446000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_932
timestamp 1765222618
transform 0 1 0 -1 0 442000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_933
timestamp 1765222618
transform 0 1 0 -1 0 438000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_934
timestamp 1765222618
transform 0 1 0 -1 0 440000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_935
timestamp 1765222618
transform 0 1 0 -1 0 436000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_936
timestamp 1765222618
transform 0 1 0 -1 0 434000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_937
timestamp 1765222618
transform 0 1 0 -1 0 430000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_938
timestamp 1765222618
transform 0 1 0 -1 0 432000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_940
timestamp 1765222618
transform 0 1 0 -1 0 405000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_941
timestamp 1765222618
transform 0 1 0 -1 0 407000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_942
timestamp 1765222618
transform 0 1 0 -1 0 413000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_943
timestamp 1765222618
transform 0 1 0 -1 0 411000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_944
timestamp 1765222618
transform 0 1 0 -1 0 409000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_945
timestamp 1765222618
transform 0 1 0 -1 0 401000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_946
timestamp 1765222618
transform 0 1 0 -1 0 403000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_947
timestamp 1765222618
transform 0 1 0 -1 0 399000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_948
timestamp 1765222618
transform 0 1 0 -1 0 397000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_949
timestamp 1765222618
transform 0 1 0 -1 0 393000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_950
timestamp 1765222618
transform 0 1 0 -1 0 395000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_951
timestamp 1765222618
transform 0 1 0 -1 0 391000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_952
timestamp 1765222618
transform 0 1 0 -1 0 389000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_955
timestamp 1765222618
transform 0 1 0 -1 0 366000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_956
timestamp 1765222618
transform 0 1 0 -1 0 368000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_957
timestamp 1765222618
transform 0 1 0 -1 0 370000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_958
timestamp 1765222618
transform 0 1 0 -1 0 362000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_959
timestamp 1765222618
transform 0 1 0 -1 0 360000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_960
timestamp 1765222618
transform 0 1 0 -1 0 364000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_961
timestamp 1765222618
transform 0 1 0 -1 0 358000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_962
timestamp 1765222618
transform 0 1 0 -1 0 354000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_963
timestamp 1765222618
transform 0 1 0 -1 0 352000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_964
timestamp 1765222618
transform 0 1 0 -1 0 356000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_965
timestamp 1765222618
transform 0 1 0 -1 0 350000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_966
timestamp 1765222618
transform 0 1 0 -1 0 348000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_967
timestamp 1765222618
transform 0 1 0 -1 0 329000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_970
timestamp 1765222618
transform 0 1 0 -1 0 325000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_971
timestamp 1765222618
transform 0 1 0 -1 0 323000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_972
timestamp 1765222618
transform 0 1 0 -1 0 327000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_973
timestamp 1765222618
transform 0 1 0 -1 0 321000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_974
timestamp 1765222618
transform 0 1 0 -1 0 317000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_975
timestamp 1765222618
transform 0 1 0 -1 0 315000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_976
timestamp 1765222618
transform 0 1 0 -1 0 319000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_977
timestamp 1765222618
transform 0 1 0 -1 0 313000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_978
timestamp 1765222618
transform 0 1 0 -1 0 309000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_979
timestamp 1765222618
transform 0 1 0 -1 0 307000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_980
timestamp 1765222618
transform 0 1 0 -1 0 311000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_981
timestamp 1765222618
transform 0 1 0 -1 0 286000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_982
timestamp 1765222618
transform 0 1 0 -1 0 288000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_985
timestamp 1765222618
transform 0 1 0 -1 0 284000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_986
timestamp 1765222618
transform 0 1 0 -1 0 272000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_987
timestamp 1765222618
transform 0 1 0 -1 0 276000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_988
timestamp 1765222618
transform 0 1 0 -1 0 274000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_989
timestamp 1765222618
transform 0 1 0 -1 0 280000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_990
timestamp 1765222618
transform 0 1 0 -1 0 278000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_991
timestamp 1765222618
transform 0 1 0 -1 0 282000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_992
timestamp 1765222618
transform 0 1 0 -1 0 270000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_993
timestamp 1765222618
transform 0 1 0 -1 0 266000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_994
timestamp 1765222618
transform 0 1 0 -1 0 268000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_995
timestamp 1765222618
transform 0 1 0 -1 0 245000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_996
timestamp 1765222618
transform 0 1 0 -1 0 247000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_999
timestamp 1765222618
transform 0 1 0 -1 0 243000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1000
timestamp 1765222618
transform 0 1 0 -1 0 231000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1001
timestamp 1765222618
transform 0 1 0 -1 0 235000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1002
timestamp 1765222618
transform 0 1 0 -1 0 233000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1003
timestamp 1765222618
transform 0 1 0 -1 0 239000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1004
timestamp 1765222618
transform 0 1 0 -1 0 237000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1005
timestamp 1765222618
transform 0 1 0 -1 0 241000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1006
timestamp 1765222618
transform 0 1 0 -1 0 227000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1007
timestamp 1765222618
transform 0 1 0 -1 0 229000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1008
timestamp 1765222618
transform 0 1 0 -1 0 225000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1009
timestamp 1765222618
transform 0 1 0 -1 0 206000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1010
timestamp 1765222618
transform 0 1 0 -1 0 204000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1011
timestamp 1765222618
transform 0 1 0 -1 0 202000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1014
timestamp 1765222618
transform 0 1 0 -1 0 200000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1015
timestamp 1765222618
transform 0 1 0 -1 0 188000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1016
timestamp 1765222618
transform 0 1 0 -1 0 190000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1017
timestamp 1765222618
transform 0 1 0 -1 0 196000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1018
timestamp 1765222618
transform 0 1 0 -1 0 198000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1019
timestamp 1765222618
transform 0 1 0 -1 0 192000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1020
timestamp 1765222618
transform 0 1 0 -1 0 194000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1021
timestamp 1765222618
transform 0 1 0 -1 0 184000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1022
timestamp 1765222618
transform 0 1 0 -1 0 186000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1025
timestamp 1765222618
transform 0 1 0 -1 0 165000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1026
timestamp 1765222618
transform 0 1 0 -1 0 163000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1027
timestamp 1765222618
transform 0 1 0 -1 0 159000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1028
timestamp 1765222618
transform 0 1 0 -1 0 161000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1029
timestamp 1765222618
transform 0 1 0 -1 0 157000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1030
timestamp 1765222618
transform 0 1 0 -1 0 155000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1031
timestamp 1765222618
transform 0 1 0 -1 0 151000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1032
timestamp 1765222618
transform 0 1 0 -1 0 153000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1033
timestamp 1765222618
transform 0 1 0 -1 0 149000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1034
timestamp 1765222618
transform 0 1 0 -1 0 147000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1035
timestamp 1765222618
transform 0 1 0 -1 0 143000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1036
timestamp 1765222618
transform 0 1 0 -1 0 145000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1038
timestamp 1765222618
transform 0 1 0 -1 0 85000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1039
timestamp 1765222618
transform 0 1 0 -1 0 83000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1040
timestamp 1765222618
transform 0 1 0 -1 0 81000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1041
timestamp 1765222618
transform 0 1 0 -1 0 79000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1042
timestamp 1765222618
transform 0 1 0 -1 0 77000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1043
timestamp 1765222618
transform 0 1 0 -1 0 73000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10  gf180mcu_ocd_io__fill10_1044
timestamp 1765222618
transform 0 1 0 -1 0 75000
box -32 13097 2032 69968
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_0
timestamp 1765303996
transform -1 0 160000 0 1 0
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_1
timestamp 1765303996
transform 1 0 230000 0 1 0
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_2
timestamp 1765303996
transform 1 0 340000 0 1 0
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_3
timestamp 1765303996
transform 1 0 395000 0 1 0
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_4
timestamp 1765303996
transform 1 0 450000 0 1 0
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_5
timestamp 1765303996
transform 1 0 505000 0 1 0
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_6
timestamp 1765303996
transform 1 0 560000 0 1 0
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_7
timestamp 1765303996
transform 0 -1 776000 1 0 104000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_8
timestamp 1765303996
transform 0 -1 776000 1 0 147000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_9
timestamp 1765303996
transform 0 -1 776000 1 0 190000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_10
timestamp 1765303996
transform 0 -1 776000 1 0 233000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_11
timestamp 1765303996
transform 0 -1 776000 1 0 276000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_12
timestamp 1765303996
transform 0 -1 776000 1 0 319000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_13
timestamp 1765303996
transform 0 -1 776000 1 0 362000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_14
timestamp 1765303996
transform 0 -1 776000 1 0 534000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_15
timestamp 1765303996
transform 0 -1 776000 1 0 577000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_16
timestamp 1765303996
transform 0 -1 776000 1 0 620000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_17
timestamp 1765303996
transform 0 -1 776000 1 0 663000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_18
timestamp 1765303996
transform 0 -1 776000 1 0 706000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_19
timestamp 1765303996
transform 0 -1 776000 1 0 749000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_20
timestamp 1765303996
transform 0 -1 776000 1 0 835000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_21
timestamp 1765303996
transform 0 -1 776000 1 0 921000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_22
timestamp 1765303996
transform -1 0 654000 0 -1 1014000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_23
timestamp 1765303996
transform -1 0 544000 0 -1 1014000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_24
timestamp 1765303996
transform -1 0 489000 0 -1 1014000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_25
timestamp 1765303996
transform -1 0 434000 0 -1 1014000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_26
timestamp 1765303996
transform -1 0 324000 0 -1 1014000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_27
timestamp 1765303996
transform -1 0 269000 0 -1 1014000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_28
timestamp 1765303996
transform -1 0 214000 0 -1 1014000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_29
timestamp 1765303996
transform -1 0 159000 0 -1 1014000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_30
timestamp 1765303996
transform -1 0 104000 0 -1 1014000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_31
timestamp 1765303996
transform 0 1 0 -1 0 905000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_32
timestamp 1765303996
transform 0 1 0 -1 0 741000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_33
timestamp 1765303996
transform 0 1 0 -1 0 700000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_34
timestamp 1765303996
transform 0 1 0 -1 0 659000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_35
timestamp 1765303996
transform 0 1 0 -1 0 618000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_36
timestamp 1765303996
transform 0 1 0 -1 0 577000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_37
timestamp 1765303996
transform 0 1 0 -1 0 536000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_38
timestamp 1765303996
transform 0 1 0 -1 0 495000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_39
timestamp 1765303996
transform 0 1 0 -1 0 372000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_40
timestamp 1765303996
transform 0 1 0 -1 0 331000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_41
timestamp 1765303996
transform 0 1 0 -1 0 290000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_42
timestamp 1765303996
transform 0 1 0 -1 0 249000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_43
timestamp 1765303996
transform 0 1 0 -1 0 208000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10x  gf180mcu_ocd_io__fill10x_44
timestamp 1765303996
transform 0 1 0 -1 0 167000
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10y  gf180mcu_ocd_io__fill10y_0
timestamp 1765303996
transform 1 0 592000 0 1 0
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10z  gf180mcu_ocd_io__fill10z_0
timestamp 1765303996
transform 1 0 507000 0 1 0
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10z  gf180mcu_ocd_io__fill10z_1
timestamp 1765303996
transform 1 0 509000 0 1 0
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10z  gf180mcu_ocd_io__fill10z_2
timestamp 1765303996
transform 1 0 511000 0 1 0
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10z  gf180mcu_ocd_io__fill10z_3
timestamp 1765303996
transform 1 0 513000 0 1 0
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10z  gf180mcu_ocd_io__fill10z_4
timestamp 1765303996
transform 1 0 515000 0 1 0
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10z  gf180mcu_ocd_io__fill10z_5
timestamp 1765303996
transform 1 0 517000 0 1 0
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10z  gf180mcu_ocd_io__fill10z_6
timestamp 1765303996
transform 1 0 519000 0 1 0
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10z  gf180mcu_ocd_io__fill10z_7
timestamp 1765303996
transform 1 0 521000 0 1 0
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10z  gf180mcu_ocd_io__fill10z_8
timestamp 1765303996
transform 1 0 523000 0 1 0
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10z  gf180mcu_ocd_io__fill10z_9
timestamp 1765303996
transform 1 0 525000 0 1 0
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10z  gf180mcu_ocd_io__fill10z_10
timestamp 1765303996
transform 1 0 527000 0 1 0
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10z  gf180mcu_ocd_io__fill10z_11
timestamp 1765303996
transform 1 0 529000 0 1 0
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10z  gf180mcu_ocd_io__fill10z_12
timestamp 1765303996
transform 1 0 531000 0 1 0
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10z  gf180mcu_ocd_io__fill10z_13
timestamp 1765303996
transform 1 0 533000 0 1 0
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10z  gf180mcu_ocd_io__fill10z_14
timestamp 1765303996
transform 1 0 535000 0 1 0
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10z  gf180mcu_ocd_io__fill10z_15
timestamp 1765303996
transform 1 0 537000 0 1 0
box -32 13097 2032 70000
use gf180mcu_ocd_io__fill10z  gf180mcu_ocd_io__fill10z_16
timestamp 1765303996
transform 1 0 590000 0 1 0
box -32 13097 2032 70000
use gf180mcu_ocd_io__bi_a  gpio_38_pad
timestamp 1765222618
transform 1 0 325000 0 1 0
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gpio_39_pad
timestamp 1765222618
transform 1 0 380000 0 1 0
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gpio_41_pad
timestamp 1765222618
transform 1 0 435000 0 1 0
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gpio_42_pad
timestamp 1765222618
transform 1 0 490000 0 1 0
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  gpio_43_pad
timestamp 1765222618
transform 1 0 545000 0 1 0
box -32 0 15032 70001
use horz_power_connect  horz_power_connect_0
timestamp 1764102312
transform 1 0 105272 0 1 70000
box 0 0 14456 200
use horz_power_connect  horz_power_connect_1
timestamp 1764102312
transform 1 0 270272 0 1 70000
box 0 0 14456 200
use horz_power_connect  horz_power_connect_2
timestamp 1764102312
transform 1 0 600272 0 1 70000
box 0 0 14456 200
use horz_power_connect  horz_power_connect_3
timestamp 1764102312
transform 1 0 655272 0 1 69999
box 0 0 14456 200
use horz_power_connect  horz_power_connect_4
timestamp 1764102312
transform 1 0 379272 0 1 943800
box 0 0 14456 200
use horz_power_connect  horz_power_connect_5
timestamp 1764102312
transform 1 0 599272 0 1 943800
box 0 0 14456 200
use gf180mcu_ocd_io__bi_a  pads[0]
timestamp 1765222618
transform 0 -1 776000 1 0 89000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[1]
timestamp 1765222618
transform 0 -1 776000 1 0 132000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[2]
timestamp 1765222618
transform 0 -1 776000 1 0 175000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[3]
timestamp 1765222618
transform 0 -1 776000 1 0 218000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[4]
timestamp 1765222618
transform 0 -1 776000 1 0 261000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[5]
timestamp 1765222618
transform 0 -1 776000 1 0 304000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[6]
timestamp 1765222618
transform 0 -1 776000 1 0 347000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[7]
timestamp 1765222618
transform 0 -1 776000 1 0 519000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[8]
timestamp 1765222618
transform 0 -1 776000 1 0 562000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[9]
timestamp 1765222618
transform 0 -1 776000 1 0 605000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[10]
timestamp 1765222618
transform 0 -1 776000 1 0 648000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[11]
timestamp 1765222618
transform 0 -1 776000 1 0 691000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[12]
timestamp 1765222618
transform 0 -1 776000 1 0 734000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[13]
timestamp 1765222618
transform 0 -1 776000 1 0 820000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[14]
timestamp 1765222618
transform 0 -1 776000 1 0 906000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[15]
timestamp 1765222618
transform -1 0 669000 0 -1 1014000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[16]
timestamp 1765222618
transform -1 0 559000 0 -1 1014000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[17]
timestamp 1765222618
transform -1 0 504000 0 -1 1014000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[18]
timestamp 1765222618
transform -1 0 449000 0 -1 1014000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[19]
timestamp 1765222618
transform -1 0 339000 0 -1 1014000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[20]
timestamp 1765222618
transform -1 0 284000 0 -1 1014000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[21]
timestamp 1765222618
transform -1 0 229000 0 -1 1014000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[22]
timestamp 1765222618
transform -1 0 174000 0 -1 1014000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[23]
timestamp 1765222618
transform -1 0 119000 0 -1 1014000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[24]
timestamp 1765222618
transform 0 1 0 -1 0 920000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[25]
timestamp 1765222618
transform 0 1 0 -1 0 756000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[26]
timestamp 1765222618
transform 0 1 0 -1 0 715000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[27]
timestamp 1765222618
transform 0 1 0 -1 0 674000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[28]
timestamp 1765222618
transform 0 1 0 -1 0 633000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[29]
timestamp 1765222618
transform 0 1 0 -1 0 592000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[30]
timestamp 1765222618
transform 0 1 0 -1 0 551000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[31]
timestamp 1765222618
transform 0 1 0 -1 0 510000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[32]
timestamp 1765222618
transform 0 1 0 -1 0 387000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[33]
timestamp 1765222618
transform 0 1 0 -1 0 346000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[34]
timestamp 1765222618
transform 0 1 0 -1 0 305000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[35]
timestamp 1765222618
transform 0 1 0 -1 0 264000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[36]
timestamp 1765222618
transform 0 1 0 -1 0 223000
box -32 0 15032 70001
use gf180mcu_ocd_io__bi_a  pads[37]
timestamp 1765222618
transform 0 1 0 -1 0 182000
box -32 0 15032 70001
use gf180mcu_ocd_io__in_s  resetb_pad $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765222618
transform 1 0 160000 0 1 0
box -32 0 15032 69970
use simple_por  simple_por_0 ../ip/simple_por/magic
timestamp 1765308861
transform 1 0 567075 0 1 1212
box 0 0 25156 8716
use gf180mcu_ocd_io__cor  user1_corner
timestamp 1765222618
transform -1 0 776000 0 -1 1014000
box 13097 13097 71000 71000
use gf180mcu_ocd_io__vdd  user1_vccd_pad $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765222618
transform 0 -1 776000 1 0 863000
box -32 0 15032 70000
use gf180mcu_ocd_io__dvdd  user1_vdda_pad_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765222618
transform 0 -1 776000 1 0 777000
box -32 0 15032 70000
use gf180mcu_ocd_io__dvdd  user1_vdda_pad_1
timestamp 1765222618
transform 0 -1 776000 1 0 476000
box -32 0 15032 70000
use gf180mcu_ocd_io__dvss  user1_vssa_pad_0 $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765222618
transform -1 0 614000 0 -1 1014000
box -32 0 15032 70000
use gf180mcu_ocd_io__dvss  user1_vssa_pad_1
timestamp 1765222618
transform 0 -1 776000 1 0 390000
box -32 0 15032 70000
use gf180mcu_ocd_io__vss  user1_vssd_pad $PDKPATH/libs.ref/gf180mcu_ocd_io/mag
timestamp 1765222618
transform 0 -1 776000 1 0 433000
box -32 0 15032 70000
use gf180mcu_ocd_io__cor  user2_corner
timestamp 1765222618
transform 1 0 0 0 -1 1014000
box 13097 13097 71000 71000
use gf180mcu_ocd_io__vdd  user2_vccd_pad
timestamp 1765222618
transform 0 1 0 -1 0 879000
box -32 0 15032 70000
use gf180mcu_ocd_io__dvdd  user2_vdda_pad
timestamp 1765222618
transform 0 1 0 -1 0 469000
box -32 0 15032 70000
use gf180mcu_ocd_io__dvss  user2_vssa_pad
timestamp 1765222618
transform 0 1 0 -1 0 797000
box -32 0 15032 70000
use gf180mcu_ocd_io__vss  user2_vssd_pad
timestamp 1765222618
transform 0 1 0 -1 0 428000
box -32 0 15032 70000
use user_id_programming  user_id_programming_0
timestamp 1764210621
transform 1 0 511654 0 -1 9172
box -86 -420 21814 1732
use gf180mcu_ocd_io__vdd  vccd_pad
timestamp 1765222618
transform 0 1 0 -1 0 100000
box -32 0 15032 70000
use gf180mcu_ocd_io__dvdd  vdda_pad
timestamp 1765222618
transform 1 0 655000 0 1 0
box -32 0 15032 70000
use gf180mcu_ocd_io__dvdd  vddio_pad_0
timestamp 1765222618
transform 0 1 0 -1 0 141000
box -32 0 15032 70000
use gf180mcu_ocd_io__dvdd  vddio_pad_1
timestamp 1765222618
transform 0 1 0 -1 0 838000
box -32 0 15032 70000
use vert_connects  vert_connects_0
timestamp 1764971740
transform 1 0 69968 0 1 166058
box 0 120 303 15270
use vert_connects  vert_connects_1
timestamp 1764971740
transform 1 0 69968 0 1 207058
box 0 120 303 15270
use vert_connects  vert_connects_2
timestamp 1764971740
transform 1 0 69968 0 1 248058
box 0 120 303 15270
use vert_connects  vert_connects_3
timestamp 1764971740
transform 1 0 69968 0 1 289058
box 0 120 303 15270
use vert_connects  vert_connects_4
timestamp 1764971740
transform 1 0 69968 0 1 330058
box 0 120 303 15270
use vert_connects  vert_connects_5
timestamp 1764971740
transform 1 0 69968 0 1 371058
box 0 120 303 15270
use vert_connects  vert_connects_6
timestamp 1764971740
transform 1 0 69968 0 1 494058
box 0 120 303 15270
use vert_connects  vert_connects_7
timestamp 1764971740
transform 1 0 69968 0 1 535058
box 0 120 303 15270
use vert_connects  vert_connects_8
timestamp 1764971740
transform 1 0 69968 0 1 576058
box 0 120 303 15270
use vert_connects  vert_connects_9
timestamp 1764971740
transform 1 0 69968 0 1 617058
box 0 120 303 15270
use vert_connects  vert_connects_10
timestamp 1764971740
transform 1 0 69968 0 1 658058
box 0 120 303 15270
use vert_connects  vert_connects_11
timestamp 1764971740
transform 1 0 69968 0 1 699058
box 0 120 303 15270
use vert_connects  vert_connects_12
timestamp 1764971740
transform 1 0 69968 0 1 740058
box 0 120 303 15270
use vert_connects  vert_connects_13
timestamp 1764971740
transform 1 0 69968 0 1 904058
box 0 120 303 15270
use vert_connects  vert_connects_14
timestamp 1764971740
transform -1 0 706032 0 -1 104942
box 0 120 303 15270
use vert_connects  vert_connects_15
timestamp 1764971740
transform -1 0 706032 0 -1 147942
box 0 120 303 15270
use vert_connects  vert_connects_16
timestamp 1764971740
transform -1 0 706032 0 -1 190942
box 0 120 303 15270
use vert_connects  vert_connects_17
timestamp 1764971740
transform -1 0 706032 0 -1 233942
box 0 120 303 15270
use vert_connects  vert_connects_18
timestamp 1764971740
transform -1 0 706032 0 -1 276942
box 0 120 303 15270
use vert_connects  vert_connects_19
timestamp 1764971740
transform -1 0 706032 0 -1 319942
box 0 120 303 15270
use vert_connects  vert_connects_20
timestamp 1764971740
transform -1 0 706032 0 -1 362942
box 0 120 303 15270
use vert_connects  vert_connects_21
timestamp 1764971740
transform -1 0 706032 0 -1 534942
box 0 120 303 15270
use vert_connects  vert_connects_22
timestamp 1764971740
transform -1 0 706032 0 -1 577942
box 0 120 303 15270
use vert_connects  vert_connects_23
timestamp 1764971740
transform -1 0 706032 0 -1 620942
box 0 120 303 15270
use vert_connects  vert_connects_24
timestamp 1764971740
transform -1 0 706032 0 -1 663942
box 0 120 303 15270
use vert_connects  vert_connects_25
timestamp 1764971740
transform -1 0 706032 0 -1 706942
box 0 120 303 15270
use vert_connects  vert_connects_26
timestamp 1764971740
transform -1 0 706032 0 -1 749942
box 0 120 303 15270
use vert_connects  vert_connects_27
timestamp 1764971740
transform -1 0 706032 0 -1 835942
box 0 120 303 15270
use vert_connects  vert_connects_28
timestamp 1764971740
transform -1 0 706032 0 -1 921942
box 0 120 303 15270
use vert_power_connect  vert_power_connect_0
timestamp 1764982451
transform 1 0 70000 0 1 85272
box 0 0 270 14456
use vert_power_connect  vert_power_connect_1
timestamp 1764982451
transform 1 0 70000 0 1 126272
box 0 0 270 14456
use vert_power_connect  vert_power_connect_2
timestamp 1764982451
transform 1 0 70000 0 1 413272
box 0 0 270 14456
use vert_power_connect  vert_power_connect_3
timestamp 1764982451
transform 1 0 70000 0 1 454272
box 0 0 270 14456
use vert_power_connect  vert_power_connect_4
timestamp 1764982451
transform 1 0 70000 0 1 782273
box 0 0 270 14456
use vert_power_connect  vert_power_connect_5
timestamp 1764982451
transform 1 0 70000 0 1 823272
box 0 0 270 14456
use vert_power_connect  vert_power_connect_6
timestamp 1764982451
transform 1 0 70000 0 1 864272
box 0 0 270 14456
use vert_power_connect  vert_power_connect_7
timestamp 1764982451
transform -1 0 706000 0 -1 404728
box 0 0 270 14456
use vert_power_connect  vert_power_connect_8
timestamp 1764982451
transform -1 0 706000 0 -1 447728
box 0 0 270 14456
use vert_power_connect  vert_power_connect_9
timestamp 1764982451
transform -1 0 706000 0 -1 490728
box 0 0 270 14456
use vert_power_connect  vert_power_connect_10
timestamp 1764982451
transform -1 0 706000 0 -1 791728
box 0 0 270 14456
use vert_power_connect  vert_power_connect_11
timestamp 1764982451
transform -1 0 706000 0 -1 877728
box 0 0 270 14456
use gf180mcu_ocd_io__dvss  vssa_pad
timestamp 1765222618
transform 1 0 105000 0 1 0
box -32 0 15032 70000
use gf180mcu_ocd_io__vss  vssd_pad
timestamp 1765222618
transform 1 0 270000 0 1 0
box -32 0 15032 70000
use gf180mcu_ocd_io__dvss  vssio_pad_0
timestamp 1765222618
transform 1 0 600000 0 1 0
box -32 0 15032 70000
use gf180mcu_ocd_io__dvss  vssio_pad_1
timestamp 1765222618
transform -1 0 394000 0 -1 1014000
box -32 0 15032 70000
<< labels >>
flabel metal2 162066 69900 162142 70200 0 FreeSans 480 90 0 0 resetb_pulldown
port 586 nsew
flabel metal2 229026 69924 229102 70200 0 FreeSans 480 90 0 0 gpio_oe[38]
port 24 nsew
flabel metal2 228880 69924 228956 70200 0 FreeSans 480 90 0 0 gpio_out[38]
port 23 nsew
flabel metal2 228734 69924 228810 70200 0 FreeSans 480 90 0 0 gpio_slew[38]
port 28 nsew
flabel metal2 217277 69924 217353 70200 0 FreeSans 480 90 0 0 gpio_ie[38]
port 22 nsew
flabel metal2 217066 69924 217142 70200 0 FreeSans 480 90 0 0 gpio_pulldown[38]
port 25 nsew
flabel metal2 216706 69923 216782 70199 0 FreeSans 480 90 0 0 gpio_ana[38]
port 490 nsew
flabel metal2 216193 69924 216269 70200 0 FreeSans 480 90 0 0 gpio_pullup[38]
port 26 nsew
flabel metal2 216564 69923 216640 70199 0 FreeSans 480 90 0 0 gpio_drive2[38]
port 20 nsew
flabel metal2 216422 69924 216498 70200 0 FreeSans 480 90 0 0 gpio_drive0[38]
port 19 nsew
flabel metal2 215672 69924 215748 70200 0 FreeSans 480 90 0 0 gpio_schmitt[38]
port 27 nsew
flabel metal2 229172 69924 229248 70200 0 FreeSans 480 90 0 0 gpio_in[38]
port 1 nsew
flabel metal2 490672 69924 490748 70200 0 FreeSans 480 90 0 0 gpio_schmitt[42]
port 625 nsew
flabel metal2 491193 69924 491269 70200 0 FreeSans 480 90 0 0 gpio_pullup[42]
port 626 nsew
flabel metal2 491422 69924 491498 70200 0 FreeSans 480 90 0 0 gpio_drive0[42]
port 627 nsew
flabel metal2 491564 69923 491640 70199 0 FreeSans 480 90 0 0 gpio_drive1[42]
port 628 nsew
flabel metal2 491706 69923 491782 70199 0 FreeSans 480 90 0 0 gpio_ana[42]
port 494 nsew
flabel metal2 492066 69924 492142 70200 0 FreeSans 480 90 0 0 gpio_pulldown[42]
port 629 nsew
flabel metal2 503734 69924 503810 70200 0 FreeSans 480 90 0 0 gpio_slew[42]
port 630 nsew
flabel metal2 435672 69924 435748 70200 0 FreeSans 480 90 0 0 gpio_schmitt[41]
port 631 nsew
flabel metal2 436193 69924 436269 70200 0 FreeSans 480 90 0 0 gpio_pullup[41]
port 632 nsew
flabel metal2 436422 69924 436498 70200 0 FreeSans 480 90 0 0 gpio_drive0[41]
port 633 nsew
flabel metal2 436564 69923 436640 70199 0 FreeSans 480 90 0 0 gpio_drive1[41]
port 634 nsew
flabel metal2 436706 69923 436782 70199 0 FreeSans 480 90 0 0 gpio_ana[41]
port 493 nsew
flabel metal2 437066 69924 437142 70200 0 FreeSans 480 90 0 0 gpio_pulldown[41]
port 635 nsew
flabel metal2 448734 69924 448810 70200 0 FreeSans 480 90 0 0 gpio_slew[41]
port 636 nsew
flabel metal2 380672 69924 380748 70200 0 FreeSans 480 90 0 0 gpio_schmitt[40]
port 637 nsew
flabel metal2 381193 69924 381269 70200 0 FreeSans 480 90 0 0 gpio_pullup[40]
port 638 nsew
flabel metal2 381422 69924 381498 70200 0 FreeSans 480 90 0 0 gpio_drive0[40]
port 639 nsew
flabel metal2 381564 69923 381640 70199 0 FreeSans 480 90 0 0 gpio_drive1[40]
port 640 nsew
flabel metal2 381706 69923 381782 70199 0 FreeSans 480 90 0 0 gpio_ana[40]
port 492 nsew
flabel metal2 382066 69924 382142 70200 0 FreeSans 480 90 0 0 gpio_pulldown[40]
port 641 nsew
flabel metal2 382277 69924 382353 70200 0 FreeSans 480 90 0 0 gpio_ie[40]
port 642 nsew
flabel metal2 393734 69924 393810 70200 0 FreeSans 480 90 0 0 gpio_slew[40]
port 643 nsew
flabel metal2 393880 69924 393956 70200 0 FreeSans 480 90 0 0 gpio_out[40]
port 644 nsew
flabel metal2 325672 69924 325748 70200 0 FreeSans 480 90 0 0 gpio_schmitt[39]
port 645 nsew
flabel metal2 326193 69924 326269 70200 0 FreeSans 480 90 0 0 gpio_pullup[39]
port 646 nsew
flabel metal2 326422 69924 326498 70200 0 FreeSans 480 90 0 0 gpio_drive0[39]
port 647 nsew
flabel metal2 326564 69923 326640 70199 0 FreeSans 480 90 0 0 gpio_drive1[39]
port 648 nsew
flabel metal2 326706 69923 326782 70199 0 FreeSans 480 90 0 0 gpio_ana[39]
port 491 nsew
flabel metal2 327066 69924 327142 70200 0 FreeSans 480 90 0 0 gpio_pulldown[39]
port 649 nsew
flabel metal2 327277 69924 327353 70200 0 FreeSans 480 90 0 0 gpio_ie[39]
port 650 nsew
flabel metal2 338734 69924 338810 70200 0 FreeSans 480 90 0 0 gpio_slew[39]
port 651 nsew
flabel metal2 338880 69924 338956 70200 0 FreeSans 480 90 0 0 gpio_out[39]
port 652 nsew
flabel metal2 339026 69924 339102 70200 0 FreeSans 480 90 0 0 gpio_oe[39]
port 7 nsew
flabel metal2 339172 69924 339248 70200 0 FreeSans 480 90 0 0 gpio_in[39]
port 6 nsew
flabel metal2 394026 69924 394102 70200 0 FreeSans 480 90 0 0 gpio_oe[40]
port 4 nsew
flabel metal2 394172 69924 394248 70200 0 FreeSans 480 90 0 0 gpio_in[40]
port 3 nsew
flabel metal2 546706 69923 546782 70199 0 FreeSans 480 90 0 0 gpio_ana[43]
port 495 nsew
flabel metal2 117218 943800 117294 944076 0 FreeSans 480 270 0 0 gpio_ana[23]
port 475 nsew
flabel metal2 172218 943800 172294 944076 0 FreeSans 480 270 0 0 gpio_ana[22]
port 474 nsew
flabel metal2 227218 943800 227294 944076 0 FreeSans 480 270 0 0 gpio_ana[21]
port 473 nsew
flabel metal2 282218 943800 282294 944076 0 FreeSans 480 270 0 0 gpio_ana[20]
port 472 nsew
flabel metal2 337218 943800 337294 944076 0 FreeSans 480 270 0 0 gpio_ana[19]
port 471 nsew
flabel metal2 447218 943800 447294 944076 0 FreeSans 480 270 0 0 gpio_ana[18]
port 470 nsew
flabel metal2 502218 943800 502294 944076 0 FreeSans 480 270 0 0 gpio_ana[17]
port 469 nsew
flabel metal2 557218 943800 557294 944076 0 FreeSans 480 270 0 0 gpio_ana[16]
port 468 nsew
flabel metal2 667218 943800 667294 944076 0 FreeSans 480 270 0 0 gpio_ana[15]
port 467 nsew
flabel metal5 400 824500 12400 836500 0 FreeSans 24000 0 0 0 vddio
port 448 nsew
flabel metal5 763600 778500 775600 790500 0 FreeSans 24000 0 0 0 vddio
port 448 nsew
flabel metal5 763600 477500 775600 489500 0 FreeSans 24000 0 0 0 vddio
port 448 nsew
flabel metal5 271500 400 283500 12400 0 FreeSans 24000 0 0 0 vssd
port 449 nsew
flabel metal5 400 414500 12400 426500 0 FreeSans 24000 0 0 0 vssd
port 449 nsew
flabel metal5 763600 434500 775600 446500 0 FreeSans 24000 0 0 0 vssd
port 449 nsew
flabel metal5 601500 400 613500 12400 0 FreeSans 24000 0 0 0 vssio
port 450 nsew
flabel metal5 106500 400 118500 12400 0 FreeSans 24000 0 0 0 vssio
port 450 nsew
flabel metal5 400 783500 12400 795500 0 FreeSans 24000 0 0 0 vssio
port 450 nsew
flabel metal5 380500 1001600 392500 1013600 0 FreeSans 24000 0 0 0 vssio
port 450 nsew
flabel metal5 600500 1001600 612500 1013600 0 FreeSans 24000 0 0 0 vssio
port 450 nsew
flabel metal5 763600 391500 775600 403500 0 FreeSans 24000 0 0 0 vssio
port 450 nsew
flabel metal5 656500 400 668500 12400 0 FreeSans 24000 0 0 0 vddio
port 448 nsew
flabel metal5 400 86500 12400 98500 0 FreeSans 24000 0 0 0 vccd
port 451 nsew
flabel metal5 400 127500 12400 139500 0 FreeSans 24000 0 0 0 vddio
port 448 nsew
flabel metal5 400 455500 12400 467500 0 FreeSans 24000 0 0 0 vddio
port 448 nsew
flabel metal5 400 865500 12400 877500 0 FreeSans 24000 0 0 0 vccd
port 451 nsew
flabel metal5 763600 864500 775600 876500 0 FreeSans 24000 0 0 0 vccd
port 451 nsew
flabel metal2 104752 943800 104828 944076 0 FreeSans 480 270 0 0 gpio_in[23]
port 157 nsew
flabel metal2 104898 943800 104974 944076 0 FreeSans 480 270 0 0 gpio_oe[23]
port 271 nsew
flabel metal2 105044 943800 105120 944076 0 FreeSans 480 270 0 0 gpio_out[23]
port 233 nsew
flabel metal2 105190 943800 105266 944076 0 FreeSans 480 270 0 0 gpio_slew[23]
port 423 nsew
flabel metal2 116647 943800 116723 944076 0 FreeSans 480 270 0 0 gpio_ie[23]
port 195 nsew
flabel metal2 116858 943800 116934 944076 0 FreeSans 480 270 0 0 gpio_pulldown[23]
port 309 nsew
flabel metal2 117360 943800 117436 944076 0 FreeSans 480 270 0 0 gpio_drive1[23]
port 108 nsew
flabel metal2 117502 943800 117578 944076 0 FreeSans 480 270 0 0 gpio_drive0[23]
port 107 nsew
flabel metal2 117731 943800 117807 944076 0 FreeSans 480 270 0 0 gpio_pullup[23]
port 347 nsew
flabel metal2 118252 943800 118328 944076 0 FreeSans 480 270 0 0 gpio_schmitt[23]
port 385 nsew
flabel metal2 159752 943800 159828 944076 0 FreeSans 480 270 0 0 gpio_in[22]
port 156 nsew
flabel metal2 159898 943800 159974 944076 0 FreeSans 480 270 0 0 gpio_oe[22]
port 270 nsew
flabel metal2 160044 943800 160120 944076 0 FreeSans 480 270 0 0 gpio_out[22]
port 232 nsew
flabel metal2 160190 943800 160266 944076 0 FreeSans 480 270 0 0 gpio_slew[22]
port 422 nsew
flabel metal2 171647 943800 171723 944076 0 FreeSans 480 270 0 0 gpio_ie[22]
port 194 nsew
flabel metal2 171858 943800 171934 944076 0 FreeSans 480 270 0 0 gpio_pulldown[22]
port 308 nsew
flabel metal2 172360 943800 172436 944076 0 FreeSans 480 270 0 0 gpio_drive1[22]
port 106 nsew
flabel metal2 172502 943800 172578 944076 0 FreeSans 480 270 0 0 gpio_drive0[22]
port 105 nsew
flabel metal2 172731 943800 172807 944076 0 FreeSans 480 270 0 0 gpio_pullup[22]
port 346 nsew
flabel metal2 173252 943800 173328 944076 0 FreeSans 480 270 0 0 gpio_schmitt[22]
port 384 nsew
flabel metal2 214752 943800 214828 944076 0 FreeSans 480 270 0 0 gpio_in[21]
port 155 nsew
flabel metal2 214898 943800 214974 944076 0 FreeSans 480 270 0 0 gpio_oe[21]
port 269 nsew
flabel metal2 215044 943800 215120 944076 0 FreeSans 480 270 0 0 gpio_out[21]
port 231 nsew
flabel metal2 215190 943800 215266 944076 0 FreeSans 480 270 0 0 gpio_slew[21]
port 421 nsew
flabel metal2 226647 943800 226723 944076 0 FreeSans 480 270 0 0 gpio_ie[21]
port 193 nsew
flabel metal2 226858 943800 226934 944076 0 FreeSans 480 270 0 0 gpio_pulldown[21]
port 307 nsew
flabel metal2 227360 943800 227436 944076 0 FreeSans 480 270 0 0 gpio_drive1[21]
port 104 nsew
flabel metal2 227502 943800 227578 944076 0 FreeSans 480 270 0 0 gpio_drive0[21]
port 103 nsew
flabel metal2 227731 943800 227807 944076 0 FreeSans 480 270 0 0 gpio_pullup[21]
port 345 nsew
flabel metal2 228252 943800 228328 944076 0 FreeSans 480 270 0 0 gpio_schmitt[21]
port 383 nsew
flabel metal2 269752 943800 269828 944076 0 FreeSans 480 270 0 0 gpio_in[20]
port 154 nsew
flabel metal2 269898 943800 269974 944076 0 FreeSans 480 270 0 0 gpio_oe[20]
port 268 nsew
flabel metal2 270044 943800 270120 944076 0 FreeSans 480 270 0 0 gpio_out[20]
port 230 nsew
flabel metal2 270190 943800 270266 944076 0 FreeSans 480 270 0 0 gpio_slew[20]
port 420 nsew
flabel metal2 281647 943800 281723 944076 0 FreeSans 480 270 0 0 gpio_ie[20]
port 192 nsew
flabel metal2 281858 943800 281934 944076 0 FreeSans 480 270 0 0 gpio_pulldown[20]
port 306 nsew
flabel metal2 282360 943800 282436 944076 0 FreeSans 480 270 0 0 gpio_drive1[20]
port 102 nsew
flabel metal2 282502 943800 282578 944076 0 FreeSans 480 270 0 0 gpio_drive0[20]
port 101 nsew
flabel metal2 282731 943800 282807 944076 0 FreeSans 480 270 0 0 gpio_pullup[20]
port 344 nsew
flabel metal2 283252 943800 283328 944076 0 FreeSans 480 270 0 0 gpio_schmitt[20]
port 382 nsew
flabel metal2 324752 943800 324828 944076 0 FreeSans 480 270 0 0 gpio_in[19]
port 152 nsew
flabel metal2 324898 943800 324974 944076 0 FreeSans 480 270 0 0 gpio_oe[19]
port 266 nsew
flabel metal2 325044 943800 325120 944076 0 FreeSans 480 270 0 0 gpio_out[19]
port 228 nsew
flabel metal2 325190 943800 325266 944076 0 FreeSans 480 270 0 0 gpio_slew[19]
port 418 nsew
flabel metal2 336647 943800 336723 944076 0 FreeSans 480 270 0 0 gpio_ie[19]
port 190 nsew
flabel metal2 336858 943800 336934 944076 0 FreeSans 480 270 0 0 gpio_pulldown[19]
port 304 nsew
flabel metal2 337360 943800 337436 944076 0 FreeSans 480 270 0 0 gpio_drive1[19]
port 99 nsew
flabel metal2 337502 943800 337578 944076 0 FreeSans 480 270 0 0 gpio_drive0[19]
port 98 nsew
flabel metal2 337731 943800 337807 944076 0 FreeSans 480 270 0 0 gpio_pullup[19]
port 342 nsew
flabel metal2 338252 943800 338328 944076 0 FreeSans 480 270 0 0 gpio_schmitt[19]
port 380 nsew
flabel metal2 434752 943800 434828 944076 0 FreeSans 480 270 0 0 gpio_in[18]
port 151 nsew
flabel metal2 434898 943800 434974 944076 0 FreeSans 480 270 0 0 gpio_oe[18]
port 265 nsew
flabel metal2 435044 943800 435120 944076 0 FreeSans 480 270 0 0 gpio_out[18]
port 227 nsew
flabel metal2 435190 943800 435266 944076 0 FreeSans 480 270 0 0 gpio_slew[18]
port 417 nsew
flabel metal2 446647 943800 446723 944076 0 FreeSans 480 270 0 0 gpio_ie[18]
port 189 nsew
flabel metal2 446858 943800 446934 944076 0 FreeSans 480 270 0 0 gpio_pulldown[18]
port 303 nsew
flabel metal2 447360 943800 447436 944076 0 FreeSans 480 270 0 0 gpio_drive1[18]
port 97 nsew
flabel metal2 447502 943800 447578 944076 0 FreeSans 480 270 0 0 gpio_drive0[18]
port 96 nsew
flabel metal2 447731 943800 447807 944076 0 FreeSans 480 270 0 0 gpio_pullup[18]
port 341 nsew
flabel metal2 448252 943800 448328 944076 0 FreeSans 480 270 0 0 gpio_schmitt[18]
port 379 nsew
flabel metal2 489752 943800 489828 944076 0 FreeSans 480 270 0 0 gpio_in[17]
port 150 nsew
flabel metal2 489898 943800 489974 944076 0 FreeSans 480 270 0 0 gpio_oe[17]
port 264 nsew
flabel metal2 490044 943800 490120 944076 0 FreeSans 480 270 0 0 gpio_out[17]
port 226 nsew
flabel metal2 490190 943800 490266 944076 0 FreeSans 480 270 0 0 gpio_slew[17]
port 416 nsew
flabel metal2 501647 943800 501723 944076 0 FreeSans 480 270 0 0 gpio_ie[17]
port 188 nsew
flabel metal2 501858 943800 501934 944076 0 FreeSans 480 270 0 0 gpio_pulldown[17]
port 302 nsew
flabel metal2 502360 943800 502436 944076 0 FreeSans 480 270 0 0 gpio_drive1[17]
port 95 nsew
flabel metal2 502502 943800 502578 944076 0 FreeSans 480 270 0 0 gpio_drive0[17]
port 94 nsew
flabel metal2 502731 943800 502807 944076 0 FreeSans 480 270 0 0 gpio_pullup[17]
port 340 nsew
flabel metal2 503252 943800 503328 944076 0 FreeSans 480 270 0 0 gpio_schmitt[17]
port 378 nsew
flabel metal2 544752 943800 544828 944076 0 FreeSans 480 270 0 0 gpio_in[16]
port 149 nsew
flabel metal2 544898 943800 544974 944076 0 FreeSans 480 270 0 0 gpio_oe[16]
port 263 nsew
flabel metal2 545044 943800 545120 944076 0 FreeSans 480 270 0 0 gpio_out[16]
port 225 nsew
flabel metal2 545190 943800 545266 944076 0 FreeSans 480 270 0 0 gpio_slew[16]
port 415 nsew
flabel metal2 556647 943800 556723 944076 0 FreeSans 480 270 0 0 gpio_ie[16]
port 187 nsew
flabel metal2 556858 943800 556934 944076 0 FreeSans 480 270 0 0 gpio_pulldown[16]
port 301 nsew
flabel metal2 557360 943800 557436 944076 0 FreeSans 480 270 0 0 gpio_drive1[16]
port 93 nsew
flabel metal2 557502 943800 557578 944076 0 FreeSans 480 270 0 0 gpio_drive0[16]
port 92 nsew
flabel metal2 557731 943800 557807 944076 0 FreeSans 480 270 0 0 gpio_pullup[16]
port 339 nsew
flabel metal2 558252 943800 558328 944076 0 FreeSans 480 270 0 0 gpio_schmitt[16]
port 377 nsew
flabel metal2 654752 943800 654828 944076 0 FreeSans 480 270 0 0 gpio_in[15]
port 148 nsew
flabel metal2 654898 943800 654974 944076 0 FreeSans 480 270 0 0 gpio_oe[15]
port 262 nsew
flabel metal2 655044 943800 655120 944076 0 FreeSans 480 270 0 0 gpio_out[15]
port 224 nsew
flabel metal2 655190 943800 655266 944076 0 FreeSans 480 270 0 0 gpio_slew[15]
port 414 nsew
flabel metal2 666647 943800 666723 944076 0 FreeSans 480 270 0 0 gpio_ie[15]
port 186 nsew
flabel metal2 666858 943800 666934 944076 0 FreeSans 480 270 0 0 gpio_pulldown[15]
port 300 nsew
flabel metal2 667360 943800 667436 944076 0 FreeSans 480 270 0 0 gpio_drive1[15]
port 91 nsew
flabel metal2 667502 943800 667578 944076 0 FreeSans 480 270 0 0 gpio_drive0[15]
port 90 nsew
flabel metal2 667731 943800 667807 944076 0 FreeSans 480 270 0 0 gpio_pullup[15]
port 338 nsew
flabel metal2 668252 943800 668328 944076 0 FreeSans 480 270 0 0 gpio_schmitt[15]
port 376 nsew
flabel metal5 105500 1001600 117500 1013600 0 FreeSans 24000 0 0 0 gpio[23]
port 44 nsew
flabel metal5 160500 1001600 172500 1013600 0 FreeSans 24000 0 0 0 gpio[22]
port 43 nsew
flabel metal5 215500 1001600 227500 1013600 0 FreeSans 24000 0 0 0 gpio[21]
port 42 nsew
flabel metal5 270500 1001600 282500 1013600 0 FreeSans 24000 0 0 0 gpio[20]
port 41 nsew
flabel metal5 325500 1001600 337500 1013600 0 FreeSans 24000 0 0 0 gpio[19]
port 39 nsew
flabel metal5 435500 1001600 447500 1013600 0 FreeSans 24000 0 0 0 gpio[18]
port 38 nsew
flabel metal5 490500 1001600 502500 1013600 0 FreeSans 24000 0 0 0 gpio[17]
port 37 nsew
flabel metal5 545500 1001600 557500 1013600 0 FreeSans 24000 0 0 0 gpio[16]
port 36 nsew
flabel metal5 655500 1001600 667500 1013600 0 FreeSans 24000 0 0 0 gpio[15]
port 35 nsew
flabel metal5 763600 907500 775600 919500 0 FreeSans 24000 0 0 0 gpio[14]
port 34 nsew
flabel metal5 763600 821500 775600 833500 0 FreeSans 24000 0 0 0 gpio[13]
port 33 nsew
flabel metal5 763600 735500 775600 747500 0 FreeSans 24000 0 0 0 gpio[12]
port 32 nsew
flabel metal5 763600 692500 775600 704500 0 FreeSans 24000 0 0 0 gpio[11]
port 31 nsew
flabel metal5 763600 649500 775600 661500 0 FreeSans 24000 0 0 0 gpio[10]
port 30 nsew
flabel metal5 763600 606500 775600 618500 0 FreeSans 24000 0 0 0 gpio[9]
port 66 nsew
flabel metal5 763600 563500 775600 575500 0 FreeSans 24000 0 0 0 gpio[8]
port 65 nsew
flabel metal5 763600 520500 775600 532500 0 FreeSans 24000 0 0 0 gpio[7]
port 64 nsew
flabel metal5 763600 348500 775600 360500 0 FreeSans 24000 0 0 0 gpio[6]
port 63 nsew
flabel metal5 763600 305500 775600 317500 0 FreeSans 24000 0 0 0 gpio[5]
port 62 nsew
flabel metal5 763600 262500 775600 274500 0 FreeSans 24000 0 0 0 gpio[4]
port 61 nsew
flabel metal5 763600 219500 775600 231500 0 FreeSans 24000 0 0 0 gpio[3]
port 60 nsew
flabel metal5 763600 176500 775600 188500 0 FreeSans 24000 0 0 0 gpio[2]
port 51 nsew
flabel metal5 763600 133500 775600 145500 0 FreeSans 24000 0 0 0 gpio[1]
port 40 nsew
flabel metal5 763600 90500 775600 102500 0 FreeSans 24000 0 0 0 gpio[0]
port 29 nsew
flabel metal5 400 168500 12400 180500 0 FreeSans 24000 0 0 0 gpio[37]
port 59 nsew
flabel metal5 400 209500 12400 221500 0 FreeSans 24000 0 0 0 gpio[36]
port 58 nsew
flabel metal5 400 250500 12400 262500 0 FreeSans 24000 0 0 0 gpio[35]
port 57 nsew
flabel metal5 400 291500 12400 303500 0 FreeSans 24000 0 0 0 gpio[34]
port 56 nsew
flabel metal5 400 332500 12400 344500 0 FreeSans 24000 0 0 0 gpio[33]
port 55 nsew
flabel metal5 400 373500 12400 385500 0 FreeSans 24000 0 0 0 gpio[32]
port 54 nsew
flabel metal5 400 496500 12400 508500 0 FreeSans 24000 0 0 0 gpio[31]
port 53 nsew
flabel metal5 400 537500 12400 549500 0 FreeSans 24000 0 0 0 gpio[30]
port 52 nsew
flabel metal5 400 578500 12400 590500 0 FreeSans 24000 0 0 0 gpio[29]
port 50 nsew
flabel metal5 400 619500 12400 631500 0 FreeSans 24000 0 0 0 gpio[28]
port 49 nsew
flabel metal5 400 660500 12400 672500 0 FreeSans 24000 0 0 0 gpio[27]
port 48 nsew
flabel metal5 400 701500 12400 713500 0 FreeSans 24000 0 0 0 gpio[26]
port 47 nsew
flabel metal5 400 742500 12400 754500 0 FreeSans 24000 0 0 0 gpio[25]
port 46 nsew
flabel metal5 400 906500 12400 918500 0 FreeSans 24000 0 0 0 gpio[24]
port 45 nsew
flabel metal2 559026 69924 559102 70200 0 FreeSans 480 90 0 0 gpio_oe[43]
port 653 nsew
flabel metal2 559172 69924 559248 70200 0 FreeSans 480 90 0 0 gpio_in[43]
port 21 nsew
flabel metal2 558880 69924 558956 70200 0 FreeSans 480 90 0 0 gpio_out[43]
port 654 nsew
flabel metal2 558734 69924 558810 70200 0 FreeSans 480 90 0 0 gpio_slew[43]
port 655 nsew
flabel metal2 547277 69924 547353 70200 0 FreeSans 480 90 0 0 gpio_ie[43]
port 656 nsew
flabel metal2 547066 69924 547142 70200 0 FreeSans 480 90 0 0 gpio_pulldown[43]
port 657 nsew
flabel metal2 546564 69923 546640 70199 0 FreeSans 480 90 0 0 gpio_drive1[43]
port 658 nsew
flabel metal2 546422 69924 546498 70200 0 FreeSans 480 90 0 0 gpio_drive0[43]
port 659 nsew
flabel metal2 546193 69924 546269 70200 0 FreeSans 480 90 0 0 gpio_pullup[43]
port 660 nsew
flabel metal2 545672 69924 545748 70200 0 FreeSans 480 90 0 0 gpio_schmitt[43]
port 661 nsew
flabel metal2 504172 69924 504248 70200 0 FreeSans 480 90 0 0 gpio_in[42]
port 14 nsew
flabel metal2 504026 69924 504102 70200 0 FreeSans 480 90 0 0 gpio_oe[42]
port 17 nsew
flabel metal2 503880 69924 503956 70200 0 FreeSans 480 90 0 0 gpio_out[42]
port 15 nsew
flabel metal2 492277 69924 492353 70200 0 FreeSans 480 90 0 0 gpio_ie[42]
port 16 nsew
flabel metal2 449171 69924 449247 70200 0 FreeSans 480 90 0 0 gpio_in[41]
port 9 nsew
flabel metal2 449026 69924 449102 70200 0 FreeSans 480 90 0 0 gpio_oe[41]
port 12 nsew
flabel metal2 448880 69924 448956 70200 0 FreeSans 480 90 0 0 gpio_out[41]
port 10 nsew
flabel metal2 437277 69924 437353 70200 0 FreeSans 480 90 0 0 gpio_ie[41]
port 11 nsew
flabel metal2 174172 69924 174248 70200 0 FreeSans 480 90 0 0 resetb_core
port 447 nsew
flabel metal5 546500 400 558500 12400 0 FreeSans 24000 0 0 0 gpio[43]
port 18 nsew
flabel metal5 491500 400 503500 12400 0 FreeSans 24000 0 0 0 gpio[42]
port 13 nsew
flabel metal5 436500 400 448500 12400 0 FreeSans 24000 0 0 0 gpio[41]
port 8 nsew
flabel metal5 381500 400 393500 12400 0 FreeSans 24000 0 0 0 gpio[40]
port 2 nsew
flabel metal5 326500 400 338500 12400 0 FreeSans 24000 0 0 0 gpio[39]
port 5 nsew
flabel metal5 161500 400 173500 12400 0 FreeSans 24000 0 0 0 resetb
port 446 nsew
flabel metal3 705730 146172 706006 146248 0 FreeSans 480 0 0 0 gpio_in[1]
port 153 nsew
flabel metal3 705730 146026 706006 146102 0 FreeSans 480 0 0 0 gpio_oe[1]
port 267 nsew
flabel metal3 705730 145880 706006 145956 0 FreeSans 480 0 0 0 gpio_out[1]
port 229 nsew
flabel metal3 705730 145734 706006 145810 0 FreeSans 480 0 0 0 gpio_slew[1]
port 419 nsew
flabel metal3 705729 133706 706005 133782 0 FreeSans 480 0 0 0 gpio_ana[1]
port 453 nsew
flabel metal3 705729 133564 706005 133640 0 FreeSans 480 0 0 0 gpio_drive1[1]
port 100 nsew
flabel metal3 705729 134277 706005 134353 0 FreeSans 480 0 0 0 gpio_ie[1]
port 191 nsew
flabel metal3 705729 134066 706005 134142 0 FreeSans 480 0 0 0 gpio_pulldown[1]
port 305 nsew
flabel metal3 705729 133422 706005 133498 0 FreeSans 480 0 0 0 gpio_drive0[1]
port 89 nsew
flabel metal3 705729 133193 706005 133269 0 FreeSans 480 0 0 0 gpio_pullup[1]
port 343 nsew
flabel metal3 705729 132672 706005 132748 0 FreeSans 480 0 0 0 gpio_schmitt[1]
port 381 nsew
flabel metal3 705729 907706 706005 907782 0 FreeSans 480 0 0 0 gpio_ana[14]
port 466 nsew
flabel metal3 705729 821706 706005 821782 0 FreeSans 480 0 0 0 gpio_ana[13]
port 465 nsew
flabel metal3 705729 735706 706005 735782 0 FreeSans 480 0 0 0 gpio_ana[12]
port 464 nsew
flabel metal3 705729 692706 706005 692782 0 FreeSans 480 0 0 0 gpio_ana[11]
port 463 nsew
flabel metal3 705729 649706 706005 649782 0 FreeSans 480 0 0 0 gpio_ana[10]
port 462 nsew
flabel metal3 705729 606706 706005 606782 0 FreeSans 480 0 0 0 gpio_ana[9]
port 461 nsew
flabel metal3 705729 563706 706005 563782 0 FreeSans 480 0 0 0 gpio_ana[8]
port 460 nsew
flabel metal3 705729 520706 706005 520782 0 FreeSans 480 0 0 0 gpio_ana[7]
port 459 nsew
flabel metal3 705729 348706 706005 348782 0 FreeSans 480 0 0 0 gpio_ana[6]
port 458 nsew
flabel metal3 705729 305706 706005 305782 0 FreeSans 480 0 0 0 gpio_ana[5]
port 457 nsew
flabel metal3 705729 262706 706005 262782 0 FreeSans 480 0 0 0 gpio_ana[4]
port 456 nsew
flabel metal3 705729 219706 706005 219782 0 FreeSans 480 0 0 0 gpio_ana[3]
port 455 nsew
flabel metal3 705729 176706 706005 176782 0 FreeSans 480 0 0 0 gpio_ana[2]
port 454 nsew
flabel metal3 705729 90706 706005 90782 0 FreeSans 480 0 0 0 gpio_ana[0]
port 452 nsew
flabel metal3 705729 735564 706005 735640 0 FreeSans 480 0 0 0 gpio_drive1[12]
port 84 nsew
flabel metal3 705729 735422 706005 735498 0 FreeSans 480 0 0 0 gpio_drive0[12]
port 83 nsew
flabel metal3 705729 692564 706005 692640 0 FreeSans 480 0 0 0 gpio_drive1[11]
port 82 nsew
flabel metal3 705729 692422 706005 692498 0 FreeSans 480 0 0 0 gpio_drive0[11]
port 81 nsew
flabel metal3 705729 649564 706005 649640 0 FreeSans 480 0 0 0 gpio_drive1[10]
port 80 nsew
flabel metal3 705729 649422 706005 649498 0 FreeSans 480 0 0 0 gpio_drive0[10]
port 79 nsew
flabel metal3 705729 606564 706005 606640 0 FreeSans 480 0 0 0 gpio_drive1[9]
port 77 nsew
flabel metal3 705729 606422 706005 606498 0 FreeSans 480 0 0 0 gpio_drive0[9]
port 76 nsew
flabel metal3 705729 563564 706005 563640 0 FreeSans 480 0 0 0 gpio_drive1[8]
port 75 nsew
flabel metal3 705729 563422 706005 563498 0 FreeSans 480 0 0 0 gpio_drive0[8]
port 74 nsew
flabel metal3 705729 520564 706005 520640 0 FreeSans 480 0 0 0 gpio_drive1[7]
port 73 nsew
flabel metal3 705729 520422 706005 520498 0 FreeSans 480 0 0 0 gpio_drive0[7]
port 72 nsew
flabel metal3 705729 348564 706005 348640 0 FreeSans 480 0 0 0 gpio_drive1[6]
port 71 nsew
flabel metal3 705729 348422 706005 348498 0 FreeSans 480 0 0 0 gpio_drive0[6]
port 70 nsew
flabel metal3 705729 305564 706005 305640 0 FreeSans 480 0 0 0 gpio_drive1[5]
port 69 nsew
flabel metal3 705729 305422 706005 305498 0 FreeSans 480 0 0 0 gpio_drive0[5]
port 68 nsew
flabel metal3 705729 262564 706005 262640 0 FreeSans 480 0 0 0 gpio_drive1[4]
port 141 nsew
flabel metal3 705729 262422 706005 262498 0 FreeSans 480 0 0 0 gpio_drive0[4]
port 140 nsew
flabel metal3 705729 219564 706005 219640 0 FreeSans 480 0 0 0 gpio_drive1[3]
port 139 nsew
flabel metal3 705729 219422 706005 219498 0 FreeSans 480 0 0 0 gpio_drive0[3]
port 132 nsew
flabel metal3 705729 176564 706005 176640 0 FreeSans 480 0 0 0 gpio_drive1[2]
port 122 nsew
flabel metal3 705729 176422 706005 176498 0 FreeSans 480 0 0 0 gpio_drive0[2]
port 111 nsew
flabel metal3 705729 820672 706005 820748 0 FreeSans 480 0 0 0 gpio_schmitt[13]
port 374 nsew
flabel metal3 705729 821193 706005 821269 0 FreeSans 480 0 0 0 gpio_pullup[13]
port 336 nsew
flabel metal3 705729 821422 706005 821498 0 FreeSans 480 0 0 0 gpio_drive0[13]
port 85 nsew
flabel metal3 705729 821564 706005 821640 0 FreeSans 480 0 0 0 gpio_drive1[13]
port 86 nsew
flabel metal3 705729 822066 706005 822142 0 FreeSans 480 0 0 0 gpio_pulldown[13]
port 298 nsew
flabel metal3 705729 822277 706005 822353 0 FreeSans 480 0 0 0 gpio_ie[13]
port 184 nsew
flabel metal3 705729 833734 706005 833810 0 FreeSans 480 0 0 0 gpio_slew[13]
port 412 nsew
flabel metal3 705729 833880 706005 833956 0 FreeSans 480 0 0 0 gpio_out[13]
port 222 nsew
flabel metal3 705729 834026 706005 834102 0 FreeSans 480 0 0 0 gpio_oe[13]
port 260 nsew
flabel metal3 705729 834172 706005 834248 0 FreeSans 480 0 0 0 gpio_in[13]
port 146 nsew
flabel metal3 705729 734672 706005 734748 0 FreeSans 480 0 0 0 gpio_schmitt[12]
port 373 nsew
flabel metal3 705729 735193 706005 735269 0 FreeSans 480 0 0 0 gpio_pullup[12]
port 335 nsew
flabel metal3 705729 736066 706005 736142 0 FreeSans 480 0 0 0 gpio_pulldown[12]
port 297 nsew
flabel metal3 705729 736277 706005 736353 0 FreeSans 480 0 0 0 gpio_ie[12]
port 183 nsew
flabel metal3 705729 747734 706005 747810 0 FreeSans 480 0 0 0 gpio_slew[12]
port 411 nsew
flabel metal3 705729 747880 706005 747956 0 FreeSans 480 0 0 0 gpio_out[12]
port 221 nsew
flabel metal3 705729 748026 706005 748102 0 FreeSans 480 0 0 0 gpio_oe[12]
port 259 nsew
flabel metal3 705729 748172 706005 748248 0 FreeSans 480 0 0 0 gpio_in[12]
port 145 nsew
flabel metal3 705729 920172 706005 920248 0 FreeSans 480 0 0 0 gpio_in[14]
port 147 nsew
flabel metal3 705729 920026 706005 920102 0 FreeSans 480 0 0 0 gpio_oe[14]
port 261 nsew
flabel metal3 705729 919880 706005 919956 0 FreeSans 480 0 0 0 gpio_out[14]
port 223 nsew
flabel metal3 705729 919734 706005 919810 0 FreeSans 480 0 0 0 gpio_slew[14]
port 413 nsew
flabel metal3 705729 908277 706005 908353 0 FreeSans 480 0 0 0 gpio_ie[14]
port 185 nsew
flabel metal3 705729 908066 706005 908142 0 FreeSans 480 0 0 0 gpio_pulldown[14]
port 299 nsew
flabel metal3 705729 907564 706005 907640 0 FreeSans 480 0 0 0 gpio_drive1[14]
port 88 nsew
flabel metal3 705729 907422 706005 907498 0 FreeSans 480 0 0 0 gpio_drive0[14]
port 87 nsew
flabel metal3 705729 907193 706005 907269 0 FreeSans 480 0 0 0 gpio_pullup[14]
port 337 nsew
flabel metal3 705729 906672 706005 906748 0 FreeSans 480 0 0 0 gpio_schmitt[14]
port 375 nsew
flabel metal3 705729 691672 706005 691748 0 FreeSans 480 0 0 0 gpio_schmitt[11]
port 372 nsew
flabel metal3 705729 692193 706005 692269 0 FreeSans 480 0 0 0 gpio_pullup[11]
port 334 nsew
flabel metal3 705729 693066 706005 693142 0 FreeSans 480 0 0 0 gpio_pulldown[11]
port 296 nsew
flabel metal3 705729 693277 706005 693353 0 FreeSans 480 0 0 0 gpio_ie[11]
port 182 nsew
flabel metal3 705729 704734 706005 704810 0 FreeSans 480 0 0 0 gpio_slew[11]
port 410 nsew
flabel metal3 705729 704880 706005 704956 0 FreeSans 480 0 0 0 gpio_out[11]
port 220 nsew
flabel metal3 705729 705026 706005 705102 0 FreeSans 480 0 0 0 gpio_oe[11]
port 258 nsew
flabel metal3 705729 705172 706005 705248 0 FreeSans 480 0 0 0 gpio_in[11]
port 144 nsew
flabel metal3 705729 648672 706005 648748 0 FreeSans 480 0 0 0 gpio_schmitt[10]
port 371 nsew
flabel metal3 705729 649193 706005 649269 0 FreeSans 480 0 0 0 gpio_pullup[10]
port 333 nsew
flabel metal3 705729 650066 706005 650142 0 FreeSans 480 0 0 0 gpio_pulldown[10]
port 295 nsew
flabel metal3 705729 650277 706005 650353 0 FreeSans 480 0 0 0 gpio_ie[10]
port 181 nsew
flabel metal3 705729 661734 706005 661810 0 FreeSans 480 0 0 0 gpio_slew[10]
port 409 nsew
flabel metal3 705729 661880 706005 661956 0 FreeSans 480 0 0 0 gpio_out[10]
port 219 nsew
flabel metal3 705729 662026 706005 662102 0 FreeSans 480 0 0 0 gpio_oe[10]
port 257 nsew
flabel metal3 705729 662172 706005 662248 0 FreeSans 480 0 0 0 gpio_in[10]
port 143 nsew
flabel metal3 705729 605672 706005 605748 0 FreeSans 480 0 0 0 gpio_schmitt[9]
port 407 nsew
flabel metal3 705729 606193 706005 606269 0 FreeSans 480 0 0 0 gpio_pullup[9]
port 369 nsew
flabel metal3 705729 607066 706005 607142 0 FreeSans 480 0 0 0 gpio_pulldown[9]
port 331 nsew
flabel metal3 705729 607277 706005 607353 0 FreeSans 480 0 0 0 gpio_ie[9]
port 217 nsew
flabel metal3 705729 618734 706005 618810 0 FreeSans 480 0 0 0 gpio_slew[9]
port 445 nsew
flabel metal3 705729 618880 706005 618956 0 FreeSans 480 0 0 0 gpio_out[9]
port 255 nsew
flabel metal3 705729 619026 706005 619102 0 FreeSans 480 0 0 0 gpio_oe[9]
port 293 nsew
flabel metal3 705729 619172 706005 619248 0 FreeSans 480 0 0 0 gpio_in[9]
port 179 nsew
flabel metal3 705729 562672 706005 562748 0 FreeSans 480 0 0 0 gpio_schmitt[8]
port 406 nsew
flabel metal3 705729 563193 706005 563269 0 FreeSans 480 0 0 0 gpio_pullup[8]
port 368 nsew
flabel metal3 705729 564066 706005 564142 0 FreeSans 480 0 0 0 gpio_pulldown[8]
port 330 nsew
flabel metal3 705729 564277 706005 564353 0 FreeSans 480 0 0 0 gpio_ie[8]
port 216 nsew
flabel metal3 705729 575734 706005 575810 0 FreeSans 480 0 0 0 gpio_slew[8]
port 444 nsew
flabel metal3 705729 575880 706005 575956 0 FreeSans 480 0 0 0 gpio_out[8]
port 254 nsew
flabel metal3 705729 576026 706005 576102 0 FreeSans 480 0 0 0 gpio_oe[8]
port 292 nsew
flabel metal3 705729 576172 706005 576248 0 FreeSans 480 0 0 0 gpio_in[8]
port 178 nsew
flabel metal3 705729 519672 706005 519748 0 FreeSans 480 0 0 0 gpio_schmitt[7]
port 405 nsew
flabel metal3 705729 520193 706005 520269 0 FreeSans 480 0 0 0 gpio_pullup[7]
port 367 nsew
flabel metal3 705729 521066 706005 521142 0 FreeSans 480 0 0 0 gpio_pulldown[7]
port 329 nsew
flabel metal3 705729 521277 706005 521353 0 FreeSans 480 0 0 0 gpio_ie[7]
port 215 nsew
flabel metal3 705729 532734 706005 532810 0 FreeSans 480 0 0 0 gpio_slew[7]
port 443 nsew
flabel metal3 705729 532880 706005 532956 0 FreeSans 480 0 0 0 gpio_out[7]
port 253 nsew
flabel metal3 705729 533026 706005 533102 0 FreeSans 480 0 0 0 gpio_oe[7]
port 291 nsew
flabel metal3 705729 533172 706005 533248 0 FreeSans 480 0 0 0 gpio_in[7]
port 177 nsew
flabel metal3 705729 347672 706005 347748 0 FreeSans 480 0 0 0 gpio_schmitt[6]
port 404 nsew
flabel metal3 705729 348193 706005 348269 0 FreeSans 480 0 0 0 gpio_pullup[6]
port 366 nsew
flabel metal3 705729 349066 706005 349142 0 FreeSans 480 0 0 0 gpio_pulldown[6]
port 328 nsew
flabel metal3 705729 349277 706005 349353 0 FreeSans 480 0 0 0 gpio_ie[6]
port 214 nsew
flabel metal3 705729 360734 706005 360810 0 FreeSans 480 0 0 0 gpio_slew[6]
port 442 nsew
flabel metal3 705729 360880 706005 360956 0 FreeSans 480 0 0 0 gpio_out[6]
port 252 nsew
flabel metal3 705729 361026 706005 361102 0 FreeSans 480 0 0 0 gpio_oe[6]
port 290 nsew
flabel metal3 705729 361172 706005 361248 0 FreeSans 480 0 0 0 gpio_in[6]
port 176 nsew
flabel metal3 705729 304672 706005 304748 0 FreeSans 480 0 0 0 gpio_schmitt[5]
port 403 nsew
flabel metal3 705729 305193 706005 305269 0 FreeSans 480 0 0 0 gpio_pullup[5]
port 365 nsew
flabel metal3 705729 306066 706005 306142 0 FreeSans 480 0 0 0 gpio_pulldown[5]
port 327 nsew
flabel metal3 705729 306277 706005 306353 0 FreeSans 480 0 0 0 gpio_ie[5]
port 213 nsew
flabel metal3 705729 317734 706005 317810 0 FreeSans 480 0 0 0 gpio_slew[5]
port 441 nsew
flabel metal3 705729 317880 706005 317956 0 FreeSans 480 0 0 0 gpio_out[5]
port 251 nsew
flabel metal3 705729 318026 706005 318102 0 FreeSans 480 0 0 0 gpio_oe[5]
port 289 nsew
flabel metal3 705729 318172 706005 318248 0 FreeSans 480 0 0 0 gpio_in[5]
port 175 nsew
flabel metal3 705729 261672 706005 261748 0 FreeSans 480 0 0 0 gpio_schmitt[4]
port 402 nsew
flabel metal3 705729 262193 706005 262269 0 FreeSans 480 0 0 0 gpio_pullup[4]
port 364 nsew
flabel metal3 705729 263066 706005 263142 0 FreeSans 480 0 0 0 gpio_pulldown[4]
port 326 nsew
flabel metal3 705729 263277 706005 263353 0 FreeSans 480 0 0 0 gpio_ie[4]
port 212 nsew
flabel metal3 705729 274734 706005 274810 0 FreeSans 480 0 0 0 gpio_slew[4]
port 440 nsew
flabel metal3 705729 274880 706005 274956 0 FreeSans 480 0 0 0 gpio_out[4]
port 250 nsew
flabel metal3 705729 275026 706005 275102 0 FreeSans 480 0 0 0 gpio_oe[4]
port 288 nsew
flabel metal3 705729 275172 706005 275248 0 FreeSans 480 0 0 0 gpio_in[4]
port 174 nsew
flabel metal3 705729 218672 706005 218748 0 FreeSans 480 0 0 0 gpio_schmitt[3]
port 401 nsew
flabel metal3 705729 219193 706005 219269 0 FreeSans 480 0 0 0 gpio_pullup[3]
port 363 nsew
flabel metal3 705729 220066 706005 220142 0 FreeSans 480 0 0 0 gpio_pulldown[3]
port 325 nsew
flabel metal3 705729 220277 706005 220353 0 FreeSans 480 0 0 0 gpio_ie[3]
port 211 nsew
flabel metal3 705729 231734 706005 231810 0 FreeSans 480 0 0 0 gpio_slew[3]
port 439 nsew
flabel metal3 705729 231880 706005 231956 0 FreeSans 480 0 0 0 gpio_out[3]
port 249 nsew
flabel metal3 705729 232026 706005 232102 0 FreeSans 480 0 0 0 gpio_oe[3]
port 287 nsew
flabel metal3 705729 232172 706005 232248 0 FreeSans 480 0 0 0 gpio_in[3]
port 173 nsew
flabel metal3 705729 175672 706005 175748 0 FreeSans 480 0 0 0 gpio_schmitt[2]
port 392 nsew
flabel metal3 705729 176193 706005 176269 0 FreeSans 480 0 0 0 gpio_pullup[2]
port 354 nsew
flabel metal3 705729 177066 706005 177142 0 FreeSans 480 0 0 0 gpio_pulldown[2]
port 316 nsew
flabel metal3 705729 177277 706005 177353 0 FreeSans 480 0 0 0 gpio_ie[2]
port 202 nsew
flabel metal3 705729 188734 706005 188810 0 FreeSans 480 0 0 0 gpio_slew[2]
port 430 nsew
flabel metal3 705729 188880 706005 188956 0 FreeSans 480 0 0 0 gpio_out[2]
port 240 nsew
flabel metal3 705729 189026 706005 189102 0 FreeSans 480 0 0 0 gpio_oe[2]
port 278 nsew
flabel metal3 705729 189172 706005 189248 0 FreeSans 480 0 0 0 gpio_in[2]
port 164 nsew
flabel metal3 705729 103172 706005 103248 0 FreeSans 480 0 0 0 gpio_in[0]
port 142 nsew
flabel metal3 705729 103026 706005 103102 0 FreeSans 480 0 0 0 gpio_oe[0]
port 256 nsew
flabel metal3 705729 102880 706005 102956 0 FreeSans 480 0 0 0 gpio_out[0]
port 218 nsew
flabel metal3 705729 102734 706005 102810 0 FreeSans 480 0 0 0 gpio_slew[0]
port 408 nsew
flabel metal3 705729 91277 706005 91353 0 FreeSans 480 0 0 0 gpio_ie[0]
port 180 nsew
flabel metal3 705729 91066 706005 91142 0 FreeSans 480 0 0 0 gpio_pulldown[0]
port 294 nsew
flabel metal3 705729 90564 706005 90640 0 FreeSans 480 0 0 0 gpio_drive1[0]
port 78 nsew
flabel metal3 705729 90422 706005 90498 0 FreeSans 480 0 0 0 gpio_drive0[0]
port 67 nsew
flabel metal3 705729 90193 706005 90269 0 FreeSans 480 0 0 0 gpio_pullup[0]
port 332 nsew
flabel metal3 705729 89672 706005 89748 0 FreeSans 480 0 0 0 gpio_schmitt[0]
port 370 nsew
flabel metal3 69995 167752 70271 167828 0 FreeSans 480 180 0 0 gpio_in[37]
port 172 nsew
flabel metal3 69995 167898 70271 167974 0 FreeSans 480 180 0 0 gpio_oe[37]
port 286 nsew
flabel metal3 69995 168044 70271 168120 0 FreeSans 480 180 0 0 gpio_out[37]
port 248 nsew
flabel metal3 69995 168190 70271 168266 0 FreeSans 480 180 0 0 gpio_slew[37]
port 438 nsew
flabel metal3 69995 179647 70271 179723 0 FreeSans 480 180 0 0 gpio_ie[37]
port 210 nsew
flabel metal3 69995 179858 70271 179934 0 FreeSans 480 180 0 0 gpio_pulldown[37]
port 324 nsew
flabel metal3 69995 180360 70271 180436 0 FreeSans 480 180 0 0 gpio_drive1[37]
port 138 nsew
flabel metal3 69995 180502 70271 180578 0 FreeSans 480 180 0 0 gpio_drive0[37]
port 137 nsew
flabel metal3 69995 180731 70271 180807 0 FreeSans 480 180 0 0 gpio_pullup[37]
port 362 nsew
flabel metal3 69995 181252 70271 181328 0 FreeSans 480 180 0 0 gpio_schmitt[37]
port 400 nsew
flabel metal3 69995 208752 70271 208828 0 FreeSans 480 180 0 0 gpio_in[36]
port 171 nsew
flabel metal3 69995 208898 70271 208974 0 FreeSans 480 180 0 0 gpio_oe[36]
port 285 nsew
flabel metal3 69995 209044 70271 209120 0 FreeSans 480 180 0 0 gpio_out[36]
port 247 nsew
flabel metal3 69995 209190 70271 209266 0 FreeSans 480 180 0 0 gpio_slew[36]
port 437 nsew
flabel metal3 69995 220647 70271 220723 0 FreeSans 480 180 0 0 gpio_ie[36]
port 209 nsew
flabel metal3 69995 220858 70271 220934 0 FreeSans 480 180 0 0 gpio_pulldown[36]
port 323 nsew
flabel metal3 69995 221360 70271 221436 0 FreeSans 480 180 0 0 gpio_drive1[36]
port 136 nsew
flabel metal3 69995 221502 70271 221578 0 FreeSans 480 180 0 0 gpio_drive0[36]
port 135 nsew
flabel metal3 69995 221731 70271 221807 0 FreeSans 480 180 0 0 gpio_pullup[36]
port 361 nsew
flabel metal3 69995 222252 70271 222328 0 FreeSans 480 180 0 0 gpio_schmitt[36]
port 399 nsew
flabel metal3 69995 249752 70271 249828 0 FreeSans 480 180 0 0 gpio_in[35]
port 170 nsew
flabel metal3 69995 249898 70271 249974 0 FreeSans 480 180 0 0 gpio_oe[35]
port 284 nsew
flabel metal3 69995 250044 70271 250120 0 FreeSans 480 180 0 0 gpio_out[35]
port 246 nsew
flabel metal3 69995 250190 70271 250266 0 FreeSans 480 180 0 0 gpio_slew[35]
port 436 nsew
flabel metal3 69995 261647 70271 261723 0 FreeSans 480 180 0 0 gpio_ie[35]
port 208 nsew
flabel metal3 69995 261858 70271 261934 0 FreeSans 480 180 0 0 gpio_pulldown[35]
port 322 nsew
flabel metal3 69995 262360 70271 262436 0 FreeSans 480 180 0 0 gpio_drive1[35]
port 134 nsew
flabel metal3 69995 262502 70271 262578 0 FreeSans 480 180 0 0 gpio_drive0[35]
port 133 nsew
flabel metal3 69995 262731 70271 262807 0 FreeSans 480 180 0 0 gpio_pullup[35]
port 360 nsew
flabel metal3 69995 263252 70271 263328 0 FreeSans 480 180 0 0 gpio_schmitt[35]
port 398 nsew
flabel metal3 69995 290752 70271 290828 0 FreeSans 480 180 0 0 gpio_in[34]
port 169 nsew
flabel metal3 69995 262218 70271 262294 0 FreeSans 480 180 0 0 gpio_ana[35]
port 487 nsew
flabel metal3 69995 221218 70271 221294 0 FreeSans 480 180 0 0 gpio_ana[36]
port 488 nsew
flabel metal3 69995 180218 70271 180294 0 FreeSans 480 180 0 0 gpio_ana[37]
port 489 nsew
flabel metal3 69995 303218 70271 303294 0 FreeSans 480 180 0 0 gpio_ana[34]
port 486 nsew
flabel metal3 69995 344218 70271 344294 0 FreeSans 480 180 0 0 gpio_ana[33]
port 485 nsew
flabel metal3 69995 385218 70271 385294 0 FreeSans 480 180 0 0 gpio_ana[32]
port 484 nsew
flabel metal3 69995 508218 70271 508294 0 FreeSans 480 180 0 0 gpio_ana[31]
port 483 nsew
flabel metal3 69995 549218 70271 549294 0 FreeSans 480 180 0 0 gpio_ana[30]
port 482 nsew
flabel metal3 69995 590218 70271 590294 0 FreeSans 480 180 0 0 gpio_ana[29]
port 481 nsew
flabel metal3 69995 631218 70271 631294 0 FreeSans 480 180 0 0 gpio_ana[28]
port 480 nsew
flabel metal3 69995 672218 70271 672294 0 FreeSans 480 180 0 0 gpio_ana[27]
port 479 nsew
flabel metal3 69995 713218 70271 713294 0 FreeSans 480 180 0 0 gpio_ana[26]
port 478 nsew
flabel metal3 69995 754218 70271 754294 0 FreeSans 480 180 0 0 gpio_ana[25]
port 477 nsew
flabel metal3 69995 918218 70271 918294 0 FreeSans 480 180 0 0 gpio_ana[24]
port 476 nsew
flabel metal3 69995 549502 70271 549578 0 FreeSans 480 180 0 0 gpio_drive0[30]
port 624 nsew
flabel metal3 69995 549360 70271 549436 0 FreeSans 480 180 0 0 gpio_drive1[30]
port 123 nsew
flabel metal3 69995 919252 70271 919328 0 FreeSans 480 180 0 0 gpio_schmitt[24]
port 386 nsew
flabel metal3 69995 918731 70271 918807 0 FreeSans 480 180 0 0 gpio_pullup[24]
port 348 nsew
flabel metal3 69995 918502 70271 918578 0 FreeSans 480 180 0 0 gpio_drive0[24]
port 109 nsew
flabel metal3 69995 918360 70271 918436 0 FreeSans 480 180 0 0 gpio_drive1[24]
port 110 nsew
flabel metal3 69995 917858 70271 917934 0 FreeSans 480 180 0 0 gpio_pulldown[24]
port 310 nsew
flabel metal3 69995 917647 70271 917723 0 FreeSans 480 180 0 0 gpio_ie[24]
port 196 nsew
flabel metal3 69995 906190 70271 906266 0 FreeSans 480 180 0 0 gpio_slew[24]
port 424 nsew
flabel metal3 69995 906044 70271 906120 0 FreeSans 480 180 0 0 gpio_out[24]
port 234 nsew
flabel metal3 69995 905898 70271 905974 0 FreeSans 480 180 0 0 gpio_oe[24]
port 272 nsew
flabel metal3 69995 905752 70271 905828 0 FreeSans 480 180 0 0 gpio_in[24]
port 158 nsew
flabel metal3 69995 755252 70271 755328 0 FreeSans 480 180 0 0 gpio_schmitt[25]
port 387 nsew
flabel metal3 69995 754731 70271 754807 0 FreeSans 480 180 0 0 gpio_pullup[25]
port 349 nsew
flabel metal3 69995 754502 70271 754578 0 FreeSans 480 180 0 0 gpio_drive0[25]
port 113 nsew
flabel metal3 69995 754360 70271 754436 0 FreeSans 480 180 0 0 gpio_drive1[25]
port 112 nsew
flabel metal3 69995 753858 70271 753934 0 FreeSans 480 180 0 0 gpio_pulldown[25]
port 311 nsew
flabel metal3 69995 753647 70271 753723 0 FreeSans 480 180 0 0 gpio_ie[25]
port 197 nsew
flabel metal3 69995 742190 70271 742266 0 FreeSans 480 180 0 0 gpio_slew[25]
port 425 nsew
flabel metal3 69995 742044 70271 742120 0 FreeSans 480 180 0 0 gpio_out[25]
port 235 nsew
flabel metal3 69995 741898 70271 741974 0 FreeSans 480 180 0 0 gpio_oe[25]
port 273 nsew
flabel metal3 69995 741752 70271 741828 0 FreeSans 480 180 0 0 gpio_in[25]
port 159 nsew
flabel metal3 69995 714252 70271 714328 0 FreeSans 480 180 0 0 gpio_schmitt[26]
port 388 nsew
flabel metal3 69995 713731 70271 713807 0 FreeSans 480 180 0 0 gpio_pullup[26]
port 350 nsew
flabel metal3 69995 713502 70271 713578 0 FreeSans 480 180 0 0 gpio_drive0[26]
port 114 nsew
flabel metal3 69995 713360 70271 713436 0 FreeSans 480 180 0 0 gpio_drive1[26]
port 115 nsew
flabel metal3 69995 712858 70271 712934 0 FreeSans 480 180 0 0 gpio_pulldown[26]
port 312 nsew
flabel metal3 69995 712647 70271 712723 0 FreeSans 480 180 0 0 gpio_ie[26]
port 198 nsew
flabel metal3 69995 701190 70271 701266 0 FreeSans 480 180 0 0 gpio_slew[26]
port 426 nsew
flabel metal3 69995 701044 70271 701120 0 FreeSans 480 180 0 0 gpio_out[26]
port 236 nsew
flabel metal3 69995 700898 70271 700974 0 FreeSans 480 180 0 0 gpio_oe[26]
port 274 nsew
flabel metal3 69995 700752 70271 700828 0 FreeSans 480 180 0 0 gpio_in[26]
port 160 nsew
flabel metal3 69995 673252 70271 673328 0 FreeSans 480 180 0 0 gpio_schmitt[27]
port 389 nsew
flabel metal3 69995 672731 70271 672807 0 FreeSans 480 180 0 0 gpio_pullup[27]
port 351 nsew
flabel metal3 69995 672502 70271 672578 0 FreeSans 480 180 0 0 gpio_drive0[27]
port 116 nsew
flabel metal3 69995 672360 70271 672436 0 FreeSans 480 180 0 0 gpio_drive1[27]
port 117 nsew
flabel metal3 69995 671858 70271 671934 0 FreeSans 480 180 0 0 gpio_pulldown[27]
port 313 nsew
flabel metal3 69995 671647 70271 671723 0 FreeSans 480 180 0 0 gpio_ie[27]
port 199 nsew
flabel metal3 69995 660190 70271 660266 0 FreeSans 480 180 0 0 gpio_slew[27]
port 427 nsew
flabel metal3 69995 660044 70271 660120 0 FreeSans 480 180 0 0 gpio_out[27]
port 237 nsew
flabel metal3 69995 659898 70271 659974 0 FreeSans 480 180 0 0 gpio_oe[27]
port 275 nsew
flabel metal3 69995 659752 70271 659828 0 FreeSans 480 180 0 0 gpio_in[27]
port 161 nsew
flabel metal3 69995 632252 70271 632328 0 FreeSans 480 180 0 0 gpio_schmitt[28]
port 390 nsew
flabel metal3 69995 631731 70271 631807 0 FreeSans 480 180 0 0 gpio_pullup[28]
port 352 nsew
flabel metal3 69995 631502 70271 631578 0 FreeSans 480 180 0 0 gpio_drive0[28]
port 118 nsew
flabel metal3 69995 631360 70271 631436 0 FreeSans 480 180 0 0 gpio_drive1[28]
port 119 nsew
flabel metal3 69995 630858 70271 630934 0 FreeSans 480 180 0 0 gpio_pulldown[28]
port 314 nsew
flabel metal3 69995 630647 70271 630723 0 FreeSans 480 180 0 0 gpio_ie[28]
port 200 nsew
flabel metal3 69995 619190 70271 619266 0 FreeSans 480 180 0 0 gpio_slew[28]
port 428 nsew
flabel metal3 69995 619044 70271 619120 0 FreeSans 480 180 0 0 gpio_out[28]
port 238 nsew
flabel metal3 69995 618898 70271 618974 0 FreeSans 480 180 0 0 gpio_oe[28]
port 276 nsew
flabel metal3 69995 618752 70271 618828 0 FreeSans 480 180 0 0 gpio_in[28]
port 162 nsew
flabel metal3 69995 591252 70271 591328 0 FreeSans 480 180 0 0 gpio_schmitt[29]
port 391 nsew
flabel metal3 69995 590731 70271 590807 0 FreeSans 480 180 0 0 gpio_pullup[29]
port 353 nsew
flabel metal3 69995 590502 70271 590578 0 FreeSans 480 180 0 0 gpio_drive0[29]
port 120 nsew
flabel metal3 69995 590360 70271 590436 0 FreeSans 480 180 0 0 gpio_drive1[29]
port 121 nsew
flabel metal3 69995 589858 70271 589934 0 FreeSans 480 180 0 0 gpio_pulldown[29]
port 315 nsew
flabel metal3 69995 589647 70271 589723 0 FreeSans 480 180 0 0 gpio_ie[29]
port 201 nsew
flabel metal3 69995 578190 70271 578266 0 FreeSans 480 180 0 0 gpio_slew[29]
port 429 nsew
flabel metal3 69995 578044 70271 578120 0 FreeSans 480 180 0 0 gpio_out[29]
port 239 nsew
flabel metal3 69995 577898 70271 577974 0 FreeSans 480 180 0 0 gpio_oe[29]
port 277 nsew
flabel metal3 69995 577752 70271 577828 0 FreeSans 480 180 0 0 gpio_in[29]
port 163 nsew
flabel metal3 69995 550252 70271 550328 0 FreeSans 480 180 0 0 gpio_schmitt[30]
port 393 nsew
flabel metal3 69995 549731 70271 549807 0 FreeSans 480 180 0 0 gpio_pullup[30]
port 355 nsew
flabel metal3 69995 548858 70271 548934 0 FreeSans 480 180 0 0 gpio_pulldown[30]
port 317 nsew
flabel metal3 69995 548647 70271 548723 0 FreeSans 480 180 0 0 gpio_ie[30]
port 203 nsew
flabel metal3 69995 537190 70271 537266 0 FreeSans 480 180 0 0 gpio_slew[30]
port 431 nsew
flabel metal3 69995 537044 70271 537120 0 FreeSans 480 180 0 0 gpio_out[30]
port 241 nsew
flabel metal3 69995 536898 70271 536974 0 FreeSans 480 180 0 0 gpio_oe[30]
port 279 nsew
flabel metal3 69995 536752 70271 536828 0 FreeSans 480 180 0 0 gpio_in[30]
port 165 nsew
flabel metal3 69995 509252 70271 509328 0 FreeSans 480 180 0 0 gpio_schmitt[31]
port 394 nsew
flabel metal3 69995 508731 70271 508807 0 FreeSans 480 180 0 0 gpio_pullup[31]
port 356 nsew
flabel metal3 69995 508502 70271 508578 0 FreeSans 480 180 0 0 gpio_drive0[31]
port 124 nsew
flabel metal3 69995 508360 70271 508436 0 FreeSans 480 180 0 0 gpio_drive1[31]
port 125 nsew
flabel metal3 69995 507858 70271 507934 0 FreeSans 480 180 0 0 gpio_pulldown[31]
port 318 nsew
flabel metal3 69995 507647 70271 507723 0 FreeSans 480 180 0 0 gpio_ie[31]
port 204 nsew
flabel metal3 69995 496190 70271 496266 0 FreeSans 480 180 0 0 gpio_slew[31]
port 432 nsew
flabel metal3 69995 496044 70271 496120 0 FreeSans 480 180 0 0 gpio_out[31]
port 242 nsew
flabel metal3 69995 495898 70271 495974 0 FreeSans 480 180 0 0 gpio_oe[31]
port 280 nsew
flabel metal3 69995 495752 70271 495828 0 FreeSans 480 180 0 0 gpio_in[31]
port 166 nsew
flabel metal3 69995 386252 70271 386328 0 FreeSans 480 180 0 0 gpio_schmitt[32]
port 395 nsew
flabel metal3 69995 385731 70271 385807 0 FreeSans 480 180 0 0 gpio_pullup[32]
port 357 nsew
flabel metal3 69995 385502 70271 385578 0 FreeSans 480 180 0 0 gpio_drive0[32]
port 126 nsew
flabel metal3 69995 385360 70271 385436 0 FreeSans 480 180 0 0 gpio_drive1[32]
port 127 nsew
flabel metal3 69995 384858 70271 384934 0 FreeSans 480 180 0 0 gpio_pulldown[32]
port 319 nsew
flabel metal3 69995 384647 70271 384723 0 FreeSans 480 180 0 0 gpio_ie[32]
port 205 nsew
flabel metal3 69995 373190 70271 373266 0 FreeSans 480 180 0 0 gpio_slew[32]
port 433 nsew
flabel metal3 69995 373044 70271 373120 0 FreeSans 480 180 0 0 gpio_out[32]
port 243 nsew
flabel metal3 69995 372898 70271 372974 0 FreeSans 480 180 0 0 gpio_oe[32]
port 281 nsew
flabel metal3 69995 372752 70271 372828 0 FreeSans 480 180 0 0 gpio_in[32]
port 167 nsew
flabel metal3 69995 345252 70271 345328 0 FreeSans 480 180 0 0 gpio_schmitt[33]
port 396 nsew
flabel metal3 69995 344731 70271 344807 0 FreeSans 480 180 0 0 gpio_pullup[33]
port 358 nsew
flabel metal3 69995 344502 70271 344578 0 FreeSans 480 180 0 0 gpio_drive0[33]
port 128 nsew
flabel metal3 69995 344360 70271 344436 0 FreeSans 480 180 0 0 gpio_drive1[33]
port 129 nsew
flabel metal3 69995 343858 70271 343934 0 FreeSans 480 180 0 0 gpio_pulldown[33]
port 320 nsew
flabel metal3 69995 343647 70271 343723 0 FreeSans 480 180 0 0 gpio_ie[33]
port 206 nsew
flabel metal3 69995 332190 70271 332266 0 FreeSans 480 180 0 0 gpio_slew[33]
port 434 nsew
flabel metal3 69995 332044 70271 332120 0 FreeSans 480 180 0 0 gpio_out[33]
port 244 nsew
flabel metal3 69995 331898 70271 331974 0 FreeSans 480 180 0 0 gpio_oe[33]
port 282 nsew
flabel metal3 69995 331752 70271 331828 0 FreeSans 480 180 0 0 gpio_in[33]
port 168 nsew
flabel metal3 69995 304252 70271 304328 0 FreeSans 480 180 0 0 gpio_schmitt[34]
port 397 nsew
flabel metal3 69995 303731 70271 303807 0 FreeSans 480 180 0 0 gpio_pullup[34]
port 359 nsew
flabel metal3 69995 303502 70271 303578 0 FreeSans 480 180 0 0 gpio_drive0[34]
port 130 nsew
flabel metal3 69995 303360 70271 303436 0 FreeSans 480 180 0 0 gpio_drive1[34]
port 131 nsew
flabel metal3 69995 302858 70271 302934 0 FreeSans 480 180 0 0 gpio_pulldown[34]
port 321 nsew
flabel metal3 69995 302647 70271 302723 0 FreeSans 480 180 0 0 gpio_ie[34]
port 207 nsew
flabel metal3 69995 291190 70271 291266 0 FreeSans 480 180 0 0 gpio_slew[34]
port 435 nsew
flabel metal3 69995 291044 70271 291120 0 FreeSans 480 180 0 0 gpio_out[34]
port 245 nsew
flabel metal3 69995 290898 70271 290974 0 FreeSans 480 180 0 0 gpio_oe[34]
port 283 nsew
flabel metal5 216500 400 228500 12400 0 FreeSans 24000 0 0 0 gpio[38]
port 0 nsew
flabel metal2 590707 69900 590783 70200 0 FreeSans 480 90 0 0 por_h
port 589 nsew
flabel metal2 593218 69900 593294 70200 0 FreeSans 480 90 0 0 porb_l
port 591 nsew
flabel metal2 508290 69900 508366 70200 0 FreeSans 480 90 0 0 mask_rev[1]
port 593 nsew
flabel metal2 511707 69900 511783 70200 0 FreeSans 480 90 0 0 mask_rev[4]
port 596 nsew
flabel metal2 512290 69900 512366 70200 0 FreeSans 480 90 0 0 mask_rev[5]
port 597 nsew
flabel metal2 513707 69900 513783 70200 0 FreeSans 480 90 0 0 mask_rev[6]
port 598 nsew
flabel metal2 514290 69900 514366 70200 0 FreeSans 480 90 0 0 mask_rev[7]
port 599 nsew
flabel metal2 515707 69900 515783 70200 0 FreeSans 480 90 0 0 mask_rev[8]
port 600 nsew
flabel metal2 516290 69900 516366 70200 0 FreeSans 480 90 0 0 mask_rev[9]
port 601 nsew
flabel metal2 517707 69900 517783 70200 0 FreeSans 480 90 0 0 mask_rev[10]
port 602 nsew
flabel metal2 518290 69900 518366 70200 0 FreeSans 480 90 0 0 mask_rev[11]
port 603 nsew
flabel metal2 519707 69900 519783 70200 0 FreeSans 480 90 0 0 mask_rev[12]
port 604 nsew
flabel metal2 520290 69900 520366 70200 0 FreeSans 480 90 0 0 mask_rev[13]
port 605 nsew
flabel metal2 521707 69900 521783 70200 0 FreeSans 480 90 0 0 mask_rev[14]
port 606 nsew
flabel metal2 522290 69900 522366 70200 0 FreeSans 480 90 0 0 mask_rev[15]
port 607 nsew
flabel metal2 523707 69900 523783 70200 0 FreeSans 480 90 0 0 mask_rev[16]
port 608 nsew
flabel metal2 524290 69900 524366 70200 0 FreeSans 480 90 0 0 mask_rev[17]
port 609 nsew
flabel metal2 525707 69900 525783 70200 0 FreeSans 480 90 0 0 mask_rev[18]
port 610 nsew
flabel metal2 526290 69900 526366 70200 0 FreeSans 480 90 0 0 mask_rev[19]
port 611 nsew
flabel metal2 527707 69900 527783 70200 0 FreeSans 480 90 0 0 mask_rev[20]
port 612 nsew
flabel metal2 528290 69900 528366 70200 0 FreeSans 480 90 0 0 mask_rev[21]
port 613 nsew
flabel metal2 529707 69900 529783 70200 0 FreeSans 480 90 0 0 mask_rev[22]
port 614 nsew
flabel metal2 530290 69900 530366 70200 0 FreeSans 480 90 0 0 mask_rev[23]
port 615 nsew
flabel metal2 531707 69900 531783 70200 0 FreeSans 480 90 0 0 mask_rev[24]
port 616 nsew
flabel metal2 532290 69900 532366 70200 0 FreeSans 480 90 0 0 mask_rev[25]
port 617 nsew
flabel metal2 533707 69900 533783 70200 0 FreeSans 480 90 0 0 mask_rev[26]
port 618 nsew
flabel metal2 534290 69900 534366 70200 0 FreeSans 480 90 0 0 mask_rev[27]
port 619 nsew
flabel metal2 535707 69900 535783 70200 0 FreeSans 480 90 0 0 mask_rev[28]
port 620 nsew
flabel metal2 536290 69900 536366 70200 0 FreeSans 480 90 0 0 mask_rev[29]
port 621 nsew
flabel metal2 537707 69900 537783 70200 0 FreeSans 480 90 0 0 mask_rev[30]
port 622 nsew
flabel metal2 538290 69900 538366 70200 0 FreeSans 480 90 0 0 mask_rev[31]
port 623 nsew
flabel metal5 70000 85272 70270 87172 0 FreeSans 1600 90 0 0 vccd
port 451 nsew
flabel metal5 70000 87752 70270 89802 0 FreeSans 1600 90 0 0 vccd
port 451 nsew
flabel metal5 70000 90122 70270 92172 0 FreeSans 1600 90 0 0 vccd
port 451 nsew
flabel metal5 70000 92828 70270 94878 0 FreeSans 1600 90 0 0 vccd
port 451 nsew
flabel metal5 70000 95198 70270 97248 0 FreeSans 1600 90 0 0 vccd
port 451 nsew
flabel metal5 70000 97828 70270 99728 0 FreeSans 1600 90 0 0 vccd
port 451 nsew
flabel metal5 70000 126272 70270 128172 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 70000 128752 70270 130802 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 70000 131122 70270 133172 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 70000 133828 70270 135878 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 70000 136198 70270 138248 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 70000 138828 70270 140728 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 70000 413272 70270 415172 0 FreeSans 1600 90 0 0 vssd
port 449 nsew
flabel metal5 70000 415752 70270 417802 0 FreeSans 1600 90 0 0 vssd
port 449 nsew
flabel metal5 70000 418122 70270 420172 0 FreeSans 1600 90 0 0 vssd
port 449 nsew
flabel metal5 70000 420828 70270 422878 0 FreeSans 1600 90 0 0 vssd
port 449 nsew
flabel metal5 70000 423198 70270 425248 0 FreeSans 1600 90 0 0 vssd
port 449 nsew
flabel metal5 70000 425828 70270 427728 0 FreeSans 1600 90 0 0 vssd
port 449 nsew
flabel metal5 70000 454272 70270 456172 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 70000 456752 70270 458802 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 70000 459122 70270 461172 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 70000 461828 70270 463878 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 70000 464198 70270 466248 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 70000 466828 70270 468728 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 70000 782273 70270 784173 0 FreeSans 1600 90 0 0 vssio
port 450 nsew
flabel metal5 70000 784753 70270 786803 0 FreeSans 1600 90 0 0 vssio
port 450 nsew
flabel metal5 70000 787123 70270 789173 0 FreeSans 1600 90 0 0 vssio
port 450 nsew
flabel metal5 70000 789829 70270 791879 0 FreeSans 1600 90 0 0 vssio
port 450 nsew
flabel metal5 70000 792199 70270 794249 0 FreeSans 1600 90 0 0 vssio
port 450 nsew
flabel metal5 70000 794829 70270 796729 0 FreeSans 1600 90 0 0 vssio
port 450 nsew
flabel metal5 70000 823272 70270 825172 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 70000 825752 70270 827802 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 70000 828122 70270 830172 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 70000 830828 70270 832878 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 70000 833198 70270 835248 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 70000 835828 70270 837728 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 70000 864272 70271 866172 0 FreeSans 1600 90 0 0 vccd
port 451 nsew
flabel metal5 70000 866752 70271 868802 0 FreeSans 1600 90 0 0 vccd
port 451 nsew
flabel metal5 70000 869122 70271 871172 0 FreeSans 1600 90 0 0 vccd
port 451 nsew
flabel metal5 70000 871828 70271 873878 0 FreeSans 1600 90 0 0 vccd
port 451 nsew
flabel metal5 70000 874198 70271 876248 0 FreeSans 1600 90 0 0 vccd
port 451 nsew
flabel metal5 70000 876828 70271 878728 0 FreeSans 1600 90 0 0 vccd
port 451 nsew
flabel metal4 379272 943800 381172 944000 0 FreeSans 1600 0 0 0 vssio
port 450 nsew
flabel metal4 381752 943800 383802 944000 0 FreeSans 1600 0 0 0 vssio
port 450 nsew
flabel metal4 384122 943800 386172 944000 0 FreeSans 1600 0 0 0 vssio
port 450 nsew
flabel metal4 386828 943800 388878 944000 0 FreeSans 1600 0 0 0 vssio
port 450 nsew
flabel metal4 389198 943800 391248 944000 0 FreeSans 1600 0 0 0 vssio
port 450 nsew
flabel metal4 391828 943800 393728 944000 0 FreeSans 1600 0 0 0 vssio
port 450 nsew
flabel metal4 599272 943800 601172 944000 0 FreeSans 1600 0 0 0 vssio
port 450 nsew
flabel metal4 601752 943800 603802 944000 0 FreeSans 1600 0 0 0 vssio
port 450 nsew
flabel metal4 604122 943800 606172 944000 0 FreeSans 1600 0 0 0 vssio
port 450 nsew
flabel metal4 606828 943800 608878 944000 0 FreeSans 1600 0 0 0 vssio
port 450 nsew
flabel metal4 609198 943800 611248 944000 0 FreeSans 1600 0 0 0 vssio
port 450 nsew
flabel metal4 611828 943800 613728 944000 0 FreeSans 1600 0 0 0 vssio
port 450 nsew
flabel metal5 705730 863272 706000 865172 0 FreeSans 1600 90 0 0 vccd
port 451 nsew
flabel metal5 705730 865752 706000 867802 0 FreeSans 1600 90 0 0 vccd
port 451 nsew
flabel metal5 705730 868122 706000 870172 0 FreeSans 1600 90 0 0 vccd
port 451 nsew
flabel metal5 705730 870828 706000 872878 0 FreeSans 1600 90 0 0 vccd
port 451 nsew
flabel metal5 705730 873198 706000 875248 0 FreeSans 1600 90 0 0 vccd
port 451 nsew
flabel metal5 705730 875828 706000 877728 0 FreeSans 1600 90 0 0 vccd
port 451 nsew
flabel metal5 705730 777272 706000 779172 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 705730 779752 706000 781802 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 705730 782122 706000 784172 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 705730 784828 706000 786878 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 705730 787198 706000 789248 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 705730 789828 706000 791728 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 705730 476272 706000 478172 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 705730 478752 706000 480802 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 705730 481122 706000 483172 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 705730 483828 706000 485878 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 705730 486198 706000 488248 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 705730 488828 706000 490728 0 FreeSans 1600 90 0 0 vddio
port 448 nsew
flabel metal5 705730 433272 706000 435172 0 FreeSans 1600 90 0 0 vssd
port 449 nsew
flabel metal5 705730 435752 706000 437802 0 FreeSans 1600 90 0 0 vssd
port 449 nsew
flabel metal5 705730 438122 706000 440172 0 FreeSans 1600 90 0 0 vssd
port 449 nsew
flabel metal5 705730 440828 706000 442878 0 FreeSans 1600 90 0 0 vssd
port 449 nsew
flabel metal5 705730 443198 706000 445248 0 FreeSans 1600 90 0 0 vssd
port 449 nsew
flabel metal5 705730 445828 706000 447728 0 FreeSans 1600 90 0 0 vssd
port 449 nsew
flabel metal5 705730 392752 706000 394802 0 FreeSans 1600 90 0 0 vssio
port 450 nsew
flabel metal5 705730 395122 706000 397172 0 FreeSans 1600 90 0 0 vssio
port 450 nsew
flabel metal5 705730 397828 706000 399878 0 FreeSans 1600 90 0 0 vssio
port 450 nsew
flabel metal5 705730 400198 706000 402248 0 FreeSans 1600 90 0 0 vssio
port 450 nsew
flabel metal5 705730 402828 706000 404728 0 FreeSans 1600 90 0 0 vssio
port 450 nsew
flabel metal4 600272 70000 602172 70200 0 FreeSans 1600 0 0 0 vssio
port 450 nsew
flabel metal4 602752 70000 604802 70200 0 FreeSans 1600 0 0 0 vssio
port 450 nsew
flabel metal4 605122 70000 607172 70200 0 FreeSans 1600 0 0 0 vssio
port 450 nsew
flabel metal4 607828 70000 609878 70200 0 FreeSans 1600 0 0 0 vssio
port 450 nsew
flabel metal4 610198 70000 612248 70200 0 FreeSans 1600 0 0 0 vssio
port 450 nsew
flabel metal4 612828 70000 614728 70200 0 FreeSans 1600 0 0 0 vssio
port 450 nsew
flabel metal4 270272 70000 272172 70200 0 FreeSans 1600 0 0 0 vssd
port 449 nsew
flabel metal4 272752 70000 274802 70200 0 FreeSans 1600 0 0 0 vssd
port 449 nsew
flabel metal4 275122 70000 277172 70200 0 FreeSans 1600 0 0 0 vssd
port 449 nsew
flabel metal4 277828 70000 279878 70200 0 FreeSans 1600 0 0 0 vssd
port 449 nsew
flabel metal4 280198 70000 282248 70200 0 FreeSans 1600 0 0 0 vssd
port 449 nsew
flabel metal4 282828 70000 284728 70200 0 FreeSans 1600 0 0 0 vssd
port 449 nsew
flabel metal4 105272 70000 107172 70200 0 FreeSans 1600 0 0 0 vssio
port 450 nsew
flabel metal4 107752 70000 109802 70200 0 FreeSans 1600 0 0 0 vssio
port 450 nsew
flabel metal4 110122 70000 112172 70200 0 FreeSans 1600 0 0 0 vssio
port 450 nsew
flabel metal4 112828 70000 114878 70200 0 FreeSans 1600 0 0 0 vssio
port 450 nsew
flabel metal4 115198 70000 117248 70200 0 FreeSans 1600 0 0 0 vssio
port 450 nsew
flabel metal4 117828 70000 119728 70200 0 FreeSans 1600 0 0 0 vssio
port 450 nsew
flabel metal4 655272 69999 657172 70199 0 FreeSans 1600 0 0 0 vddio
port 448 nsew
flabel metal4 657752 69999 659802 70199 0 FreeSans 1600 0 0 0 vddio
port 448 nsew
flabel metal4 660122 69999 662172 70199 0 FreeSans 1600 0 0 0 vddio
port 448 nsew
flabel metal4 662828 69999 664878 70199 0 FreeSans 1600 0 0 0 vddio
port 448 nsew
flabel metal4 665198 69999 667248 70199 0 FreeSans 1600 0 0 0 vddio
port 448 nsew
flabel metal4 667828 69999 669728 70199 0 FreeSans 1600 0 0 0 vddio
port 448 nsew
flabel metal3 705729 104746 706029 104822 0 FreeSans 480 0 0 0 gpio_loopback_zero[0]
port 496 nsew
flabel metal3 705729 104558 706029 104634 0 FreeSans 480 0 0 0 gpio_loopback_one[0]
port 497 nsew
flabel metal3 705729 147746 706029 147822 0 FreeSans 480 0 0 0 gpio_loopback_zero[1]
port 498 nsew
flabel metal3 705729 147558 706029 147634 0 FreeSans 480 0 0 0 gpio_loopback_one[1]
port 499 nsew
flabel metal3 705729 190746 706029 190822 0 FreeSans 480 0 0 0 gpio_loopback_zero[2]
port 500 nsew
flabel metal3 705729 190558 706029 190634 0 FreeSans 480 0 0 0 gpio_loopback_one[2]
port 501 nsew
flabel metal3 705729 233558 706029 233634 0 FreeSans 480 0 0 0 gpio_loopback_one[3]
port 502 nsew
flabel metal3 705729 233746 706029 233822 0 FreeSans 480 0 0 0 gpio_loopback_zero[3]
port 503 nsew
flabel metal3 705729 276558 706029 276634 0 FreeSans 480 0 0 0 gpio_loopback_one[4]
port 505 nsew
flabel metal3 705729 276746 706029 276822 0 FreeSans 480 0 0 0 gpio_loopback_zero[4]
port 504 nsew
flabel metal3 705729 319558 706029 319634 0 FreeSans 480 0 0 0 gpio_loopback_one[5]
port 506 nsew
flabel metal3 705729 319746 706029 319822 0 FreeSans 480 0 0 0 gpio_loopback_zero[5]
port 507 nsew
flabel metal3 705729 362558 706029 362634 0 FreeSans 480 0 0 0 gpio_loopback_one[6]
port 509 nsew
flabel metal3 705729 362746 706029 362822 0 FreeSans 480 0 0 0 gpio_loopback_zero[6]
port 508 nsew
flabel metal3 705729 534558 706029 534634 0 FreeSans 480 0 0 0 gpio_loopback_one[7]
port 510 nsew
flabel metal3 705729 534746 706029 534822 0 FreeSans 480 0 0 0 gpio_loopback_zero[7]
port 511 nsew
flabel metal3 705729 577558 706029 577634 0 FreeSans 480 0 0 0 gpio_loopback_one[8]
port 513 nsew
flabel metal3 705729 577746 706029 577822 0 FreeSans 480 0 0 0 gpio_loopback_zero[8]
port 512 nsew
flabel metal3 705729 620558 706029 620634 0 FreeSans 480 0 0 0 gpio_loopback_one[9]
port 514 nsew
flabel metal3 705729 620746 706029 620822 0 FreeSans 480 0 0 0 gpio_loopback_zero[9]
port 515 nsew
flabel metal3 705729 663558 706029 663634 0 FreeSans 480 0 0 0 gpio_loopback_one[10]
port 517 nsew
flabel metal3 705729 663746 706029 663822 0 FreeSans 480 0 0 0 gpio_loopback_zero[10]
port 516 nsew
flabel metal3 705729 749558 706029 749634 0 FreeSans 480 0 0 0 gpio_loopback_one[12]
port 521 nsew
flabel metal3 705729 749746 706029 749822 0 FreeSans 480 0 0 0 gpio_loopback_zero[12]
port 520 nsew
flabel metal3 705729 835558 706029 835634 0 FreeSans 480 0 0 0 gpio_loopback_one[13]
port 522 nsew
flabel metal3 705729 835746 706029 835822 0 FreeSans 480 0 0 0 gpio_loopback_zero[13]
port 523 nsew
flabel metal3 705729 921558 706029 921634 0 FreeSans 480 0 0 0 gpio_loopback_one[14]
port 525 nsew
flabel metal3 705729 921746 706029 921822 0 FreeSans 480 0 0 0 gpio_loopback_zero[14]
port 524 nsew
flabel metal2 653178 943800 653254 944100 0 FreeSans 480 90 0 0 gpio_loopback_zero[15]
port 527 nsew
flabel metal2 653366 943800 653442 944100 0 FreeSans 480 90 0 0 gpio_loopback_one[15]
port 526 nsew
flabel metal2 543366 943800 543422 944100 0 FreeSans 480 90 0 0 gpio_loopback_one[16]
port 529 nsew
flabel metal2 543178 943800 543254 944100 0 FreeSans 480 90 0 0 gpio_loopback_zero[16]
port 528 nsew
flabel metal2 488366 943800 488442 944100 0 FreeSans 480 90 0 0 gpio_loopback_one[17]
port 530 nsew
flabel metal2 488178 943800 488254 944100 0 FreeSans 480 90 0 0 gpio_loopback_zero[17]
port 531 nsew
flabel metal2 433366 943800 433442 944100 0 FreeSans 480 90 0 0 gpio_loopback_one[18]
port 533 nsew
flabel metal2 433178 943800 433254 944100 0 FreeSans 480 90 0 0 gpio_loopback_zero[18]
port 532 nsew
flabel metal2 323366 943800 323442 944100 0 FreeSans 480 90 0 0 gpio_loopback_one[19]
port 534 nsew
flabel metal2 323178 943800 323254 944100 0 FreeSans 480 90 0 0 gpio_loopback_zero[19]
port 535 nsew
flabel metal2 268366 943800 268442 944100 0 FreeSans 480 90 0 0 gpio_loopback_one[20]
port 537 nsew
flabel metal2 268178 943800 268254 944100 0 FreeSans 480 90 0 0 gpio_loopback_zero[20]
port 536 nsew
flabel metal2 213366 943800 213442 944100 0 FreeSans 480 90 0 0 gpio_loopback_one[21]
port 538 nsew
flabel metal2 213178 943800 213254 944100 0 FreeSans 480 90 0 0 gpio_loopback_zero[21]
port 539 nsew
flabel metal2 158366 943800 158442 944100 0 FreeSans 480 90 0 0 gpio_loopback_one[22]
port 541 nsew
flabel metal2 158178 943800 158254 944100 0 FreeSans 480 90 0 0 gpio_loopback_zero[22]
port 540 nsew
flabel metal2 103366 943800 103442 944100 0 FreeSans 480 90 0 0 gpio_loopback_one[23]
port 542 nsew
flabel metal2 103178 943800 103254 944100 0 FreeSans 480 90 0 0 gpio_loopback_zero[23]
port 543 nsew
flabel metal3 69971 904366 70271 904442 0 FreeSans 480 0 0 0 gpio_loopback_one[24]
port 545 nsew
flabel metal3 69971 904178 70271 904254 0 FreeSans 480 0 0 0 gpio_loopback_zero[24]
port 544 nsew
flabel metal3 69971 740366 70271 740442 0 FreeSans 480 0 0 0 gpio_loopback_one[25]
port 546 nsew
flabel metal3 69971 740178 70271 740254 0 FreeSans 480 0 0 0 gpio_loopback_zero[25]
port 547 nsew
flabel metal3 69971 699366 70271 699442 0 FreeSans 480 0 0 0 gpio_loopback_one[26]
port 549 nsew
flabel metal3 69971 699178 70271 699254 0 FreeSans 480 0 0 0 gpio_loopback_zero[26]
port 548 nsew
flabel metal3 69971 658366 70271 658442 0 FreeSans 480 0 0 0 gpio_loopback_one[27]
port 550 nsew
flabel metal3 69971 658178 70271 658254 0 FreeSans 480 0 0 0 gpio_loopback_zero[27]
port 551 nsew
flabel metal3 69971 617366 70271 617442 0 FreeSans 480 0 0 0 gpio_loopback_one[28]
port 553 nsew
flabel metal3 69971 617178 70271 617254 0 FreeSans 480 0 0 0 gpio_loopback_zero[28]
port 552 nsew
flabel metal3 69971 576366 70271 576442 0 FreeSans 480 0 0 0 gpio_loopback_one[29]
port 554 nsew
flabel metal3 69971 576178 70271 576254 0 FreeSans 480 0 0 0 gpio_loopback_zero[29]
port 555 nsew
flabel metal3 69971 535366 70271 535442 0 FreeSans 480 0 0 0 gpio_loopback_one[30]
port 557 nsew
flabel metal3 69971 535178 70271 535254 0 FreeSans 480 0 0 0 gpio_loopback_zero[30]
port 556 nsew
flabel metal3 69971 494366 70271 494442 0 FreeSans 480 0 0 0 gpio_loopback_one[31]
port 558 nsew
flabel metal3 69971 494178 70271 494254 0 FreeSans 480 0 0 0 gpio_loopback_zero[31]
port 559 nsew
flabel metal3 69971 371366 70271 371442 0 FreeSans 480 0 0 0 gpio_loopback_one[32]
port 561 nsew
flabel metal3 69971 371178 70271 371254 0 FreeSans 480 0 0 0 gpio_loopback_zero[32]
port 560 nsew
flabel metal3 69971 330366 70271 330442 0 FreeSans 480 0 0 0 gpio_loopback_one[33]
port 562 nsew
flabel metal3 69971 330178 70271 330254 0 FreeSans 480 0 0 0 gpio_loopback_zero[33]
port 563 nsew
flabel metal3 69971 289366 70271 289442 0 FreeSans 480 0 0 0 gpio_loopback_one[34]
port 565 nsew
flabel metal3 69971 289178 70271 289254 0 FreeSans 480 0 0 0 gpio_loopback_zero[34]
port 564 nsew
flabel metal3 69971 248366 70271 248442 0 FreeSans 480 0 0 0 gpio_loopback_one[35]
port 566 nsew
flabel metal3 69971 248178 70271 248254 0 FreeSans 480 0 0 0 gpio_loopback_zero[35]
port 567 nsew
flabel metal3 69971 207366 70271 207442 0 FreeSans 480 0 0 0 gpio_loopback_one[36]
port 569 nsew
flabel metal3 69971 207178 70271 207254 0 FreeSans 480 0 0 0 gpio_loopback_zero[36]
port 568 nsew
flabel metal3 69971 166366 70271 166442 0 FreeSans 480 0 0 0 gpio_loopback_one[37]
port 570 nsew
flabel metal3 69971 166178 70271 166254 0 FreeSans 480 0 0 0 gpio_loopback_zero[37]
port 571 nsew
flabel metal2 159366 69900 159442 70200 0 FreeSans 480 90 0 0 resetb_loopback_one
port 587 nsew
flabel metal2 159178 69900 159254 70200 0 FreeSans 480 90 0 0 resetb_loopback_zero
port 588 nsew
flabel metal2 230746 69900 230822 70200 0 FreeSans 480 90 0 0 gpio_loopback_zero[38]
port 572 nsew
flabel metal2 230558 69900 230634 70200 0 FreeSans 480 90 0 0 gpio_loopback_one[38]
port 573 nsew
flabel metal2 340558 69900 340634 70200 0 FreeSans 480 90 0 0 gpio_loopback_one[39]
port 574 nsew
flabel metal2 340746 69900 340822 70200 0 FreeSans 480 90 0 0 gpio_loopback_zero[39]
port 576 nsew
flabel metal2 395558 69900 395634 70200 0 FreeSans 480 90 0 0 gpio_loopback_one[40]
port 578 nsew
flabel metal2 395746 69900 395822 70200 0 FreeSans 480 90 0 0 gpio_loopback_zero[40]
port 577 nsew
flabel metal2 450558 69900 450634 70200 0 FreeSans 480 90 0 0 gpio_loopback_one[41]
port 579 nsew
flabel metal2 450746 69900 450822 70200 0 FreeSans 480 90 0 0 gpio_loopback_zero[41]
port 580 nsew
flabel metal2 505558 69900 505634 70200 0 FreeSans 480 90 0 0 gpio_loopback_one[42]
port 582 nsew
flabel metal2 505746 69900 505822 70200 0 FreeSans 480 90 0 0 gpio_loopback_zero[42]
port 581 nsew
flabel metal2 560558 69900 560634 70200 0 FreeSans 480 90 0 0 gpio_loopback_one[43]
port 583 nsew
flabel metal2 560746 69900 560822 70200 0 FreeSans 480 90 0 0 gpio_loopback_zero[43]
port 584 nsew
flabel metal3 705729 706746 706029 706822 0 FreeSans 480 0 0 0 gpio_loopback_zero[11]
port 519 nsew
flabel metal3 705729 706558 706029 706634 0 FreeSans 480 0 0 0 gpio_loopback_one[11]
port 518 nsew
flabel metal5 705730 390272 706000 392172 0 FreeSans 1600 90 0 0 vssio
port 450 nsew
flabel metal2 161194 69900 161270 70200 0 FreeSans 480 90 0 0 resetb_pullup
port 585 nsew
flabel metal2 507707 69900 507783 70200 0 FreeSans 480 90 0 0 mask_rev[0]
port 592 nsew
flabel metal2 591290 69900 591366 70200 0 FreeSans 480 90 0 0 porb_h
port 590 nsew
flabel metal2 510290 69900 510366 70200 0 FreeSans 480 90 0 0 mask_rev[3]
port 595 nsew
flabel metal2 509707 69900 509783 70200 0 FreeSans 480 90 0 0 mask_rev[2]
port 594 nsew
<< end >>
