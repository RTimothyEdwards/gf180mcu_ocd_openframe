magic
tech gf180mcuD
magscale 1 10
timestamp 1765307558
<< checkpaint >>
rect -2000 -2000 788400 1026400
<< psubdiff >>
tri 0 1022600 1800 1024400 se
rect 1800 1022600 784600 1024400
tri 784600 1022600 786400 1024400 sw
rect 0 1021200 786400 1022600
rect 0 3200 3200 1021200
rect 783200 3200 786400 1021200
rect 0 1800 786400 3200
tri 0 0 1800 1800 ne
rect 1800 0 784600 1800
tri 784600 0 786400 1800 nw
<< metal1 >>
tri 939 1023539 1800 1024400 se
rect 1800 1023539 784600 1024400
tri 665 1023265 939 1023539 se
rect 939 1023265 784600 1023539
tri 619 1023219 665 1023265 se
rect 665 1023219 784600 1023265
tri 299 1022899 619 1023219 se
rect 619 1022899 784600 1023219
tri 0 1022600 299 1022899 se
rect 299 1022600 784600 1022899
tri 784600 1022600 786400 1024400 sw
rect 0 1021400 786400 1022600
rect 0 3000 3000 1021400
tri 3000 1021200 3200 1021400 nw
tri 783200 1021200 783400 1021400 ne
tri 3000 3000 3200 3200 sw
tri 783200 3000 783400 3200 se
rect 783400 3000 786400 1021400
rect 0 1800 786400 3000
tri 0 0 1800 1800 ne
rect 1800 0 784600 1800
tri 784600 0 786400 1800 nw
<< metal2 >>
tri 1288 1023888 1800 1024400 se
rect 1800 1023888 784600 1024400
tri 928 1023528 1288 1023888 se
rect 1288 1023528 784600 1023888
tri 568 1023168 928 1023528 se
rect 928 1023168 784600 1023528
tri 0 1022600 568 1023168 se
rect 568 1022600 784600 1023168
tri 784600 1022600 786400 1024400 sw
rect 0 1021200 786400 1022600
rect 0 3200 3200 1021200
rect 783200 3200 786400 1021200
rect 0 1800 786400 3200
tri 0 0 1800 1800 ne
rect 1800 0 784600 1800
tri 784600 0 786400 1800 nw
<< metal3 >>
tri 0 1022600 1800 1024400 se
rect 1800 1022600 784600 1024400
tri 784600 1022600 786400 1024400 sw
rect 0 1021400 786400 1022600
rect 0 3000 3000 1021400
tri 3000 1021200 3200 1021400 nw
tri 783200 1021200 783400 1021400 ne
tri 3000 3000 3200 3200 sw
tri 783200 3000 783400 3200 se
rect 783400 3000 786400 1021400
rect 0 1800 786400 3000
tri 0 0 1800 1800 ne
rect 1800 0 784600 1800
tri 784600 0 786400 1800 nw
<< metal4 >>
tri 0 1022600 1800 1024400 se
rect 1800 1022600 784600 1024400
tri 784600 1022600 786400 1024400 sw
rect 0 1021200 786400 1022600
rect 0 3200 3200 1021200
rect 783200 3200 786400 1021200
rect 0 1800 786400 3200
tri 0 0 1800 1800 ne
rect 1800 0 784600 1800
tri 784600 0 786400 1800 nw
<< metal5 >>
tri 0 1022600 1800 1024400 se
rect 1800 1022600 784600 1024400
tri 784600 1022600 786400 1024400 sw
rect 0 1021400 786400 1022600
rect 0 3000 3000 1021400
tri 3000 1021200 3200 1021400 nw
tri 783200 1021200 783400 1021400 ne
tri 3000 3000 3200 3200 sw
tri 783200 3000 783400 3200 se
rect 783400 3000 786400 1021400
rect 0 1800 786400 3000
tri 0 0 1800 1800 ne
rect 1800 0 784600 1800
tri 784600 0 786400 1800 nw
<< glass >>
tri 600 1022000 2400 1023800 se
rect 2400 1022000 784000 1023800
tri 784000 1022000 785800 1023800 sw
rect 600 2400 2400 1022000
tri 2400 1021200 3200 1022000 nw
tri 783200 1021200 784000 1022000 ne
tri 2400 2400 3200 3200 sw
tri 783200 2400 784000 3200 se
rect 784000 2400 785800 1022000
tri 600 600 2400 2400 ne
rect 2400 600 784000 2400
tri 784000 600 785800 2400 nw
<< properties >>
string GDS_END 39917948
string GDS_FILE ../gds/wafer_space_sealring.gds.gz
string GDS_START 104
<< end >>
