magic
tech gf180mcuD
magscale 1 10
timestamp 1764170366
<< metal1 >>
rect 0 133 14910 185
rect 15076 133 15452 185
rect 0 35 15270 87
rect 15436 35 15452 87
<< via1 >>
rect 14910 133 15076 185
rect 15270 35 15436 87
<< metal2 >>
rect 182 0 258 232
rect 703 0 779 232
rect 932 0 1008 232
rect 1074 0 1150 232
rect 1216 0 1292 232
rect 1576 0 1652 232
rect 1787 0 1863 232
rect 13244 0 13320 232
rect 13390 0 13466 232
rect 13536 0 13612 232
rect 13682 0 13758 232
rect 15089 187 15145 232
rect 14898 185 15145 187
rect 14898 133 14910 185
rect 15076 133 15145 185
rect 14898 131 15145 133
rect 15089 0 15145 131
rect 15201 89 15257 232
rect 15201 87 15448 89
rect 15201 35 15270 87
rect 15436 35 15448 87
rect 15201 33 15448 35
rect 15201 0 15257 33
<< end >>
