magic
tech gf180mcuD
magscale 1 10
timestamp 1765308861
<< metal1 >>
rect -41 -212 2 -160
rect 54 -212 97 -160
<< via1 >>
rect 2 -212 54 -160
<< metal2 >>
rect -43 -160 99 -158
rect -43 -212 2 -160
rect 54 -212 99 -160
rect -43 -214 99 -212
<< properties >>
string GDS_END 80098
string GDS_FILE ../gds/simple_por.gds.gz
string GDS_START 79902
<< end >>
