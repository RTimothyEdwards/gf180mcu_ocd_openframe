magic
tech gf180mcuD
magscale 1 10
timestamp 1764985423
<< via1 >>
rect 161206 70101 161258 70153
rect 162079 70003 162131 70055
<< metal2 >>
rect 103178 943800 103254 944188
rect 103366 943800 103442 944188
rect 104752 943800 104828 944188
rect 104898 943800 104974 944188
rect 105044 943800 105120 944188
rect 105190 943800 105266 944188
rect 116647 943800 116723 944188
rect 116858 943800 116934 944188
rect 117218 943800 117294 944188
rect 117360 943800 117436 944188
rect 117502 943800 117578 944188
rect 117731 943800 117807 944188
rect 118252 943800 118328 944188
rect 158178 943800 158254 944188
rect 158366 943800 158442 944188
rect 159752 943800 159828 944188
rect 159898 943800 159974 944188
rect 160044 943800 160120 944188
rect 160190 943800 160266 944188
rect 171647 943800 171723 944188
rect 171858 943800 171934 944188
rect 172218 943800 172294 944188
rect 172360 943800 172436 944188
rect 172502 943800 172578 944188
rect 172731 943800 172807 944188
rect 173252 943800 173328 944188
rect 213178 943800 213254 944188
rect 213366 943800 213442 944188
rect 214752 943800 214828 944188
rect 214898 943800 214974 944188
rect 215044 943800 215120 944188
rect 215190 943800 215266 944188
rect 226647 943800 226723 944188
rect 226858 943800 226934 944188
rect 227218 943800 227294 944188
rect 227360 943800 227436 944188
rect 227502 943800 227578 944188
rect 227731 943800 227807 944188
rect 228252 943800 228328 944188
rect 268178 943800 268254 944188
rect 268366 943800 268442 944188
rect 269752 943800 269828 944188
rect 269898 943800 269974 944188
rect 270044 943800 270120 944188
rect 270190 943800 270266 944188
rect 281647 943800 281723 944188
rect 281858 943800 281934 944188
rect 282218 943800 282294 944188
rect 282360 943800 282436 944188
rect 282502 943800 282578 944188
rect 282731 943800 282807 944188
rect 283252 943800 283328 944188
rect 323178 943800 323254 944188
rect 323366 943800 323442 944188
rect 324752 943800 324828 944188
rect 324898 943800 324974 944188
rect 325044 943800 325120 944188
rect 325190 943800 325266 944188
rect 336647 943800 336723 944188
rect 336858 943800 336934 944188
rect 337218 943800 337294 944188
rect 337360 943800 337436 944188
rect 337502 943800 337578 944188
rect 337731 943800 337807 944188
rect 338252 943800 338328 944188
rect 433178 943800 433254 944188
rect 433366 943800 433442 944188
rect 434752 943800 434828 944188
rect 434898 943800 434974 944188
rect 435044 943800 435120 944188
rect 435190 943800 435266 944188
rect 446647 943800 446723 944188
rect 446858 943800 446934 944188
rect 447218 943800 447294 944188
rect 447360 943800 447436 944188
rect 447502 943800 447578 944188
rect 447731 943800 447807 944188
rect 448252 943800 448328 944188
rect 488178 943800 488254 944188
rect 488366 943800 488442 944188
rect 489752 943800 489828 944188
rect 489898 943800 489974 944188
rect 490044 943800 490120 944188
rect 490190 943800 490266 944188
rect 501647 943800 501723 944188
rect 501858 943800 501934 944188
rect 502218 943800 502294 944188
rect 502360 943800 502436 944188
rect 502502 943800 502578 944188
rect 502731 943800 502807 944188
rect 503252 943800 503328 944188
rect 543178 943800 543254 944188
rect 543366 943800 543442 944188
rect 544752 943800 544828 944188
rect 544898 943800 544974 944188
rect 545044 943800 545120 944188
rect 545190 943800 545266 944188
rect 556647 943800 556723 944188
rect 556858 943800 556934 944188
rect 557218 943800 557294 944188
rect 557360 943800 557436 944188
rect 557502 943800 557578 944188
rect 557731 943800 557807 944188
rect 558252 943800 558328 944188
rect 653178 943800 653254 944188
rect 653366 943800 653442 944188
rect 654752 943800 654828 944188
rect 654898 943800 654974 944188
rect 655044 943800 655120 944188
rect 655190 943800 655266 944188
rect 666647 943800 666723 944188
rect 666858 943800 666934 944188
rect 667218 943800 667294 944188
rect 667360 943800 667436 944188
rect 667502 943800 667578 944188
rect 667731 943800 667807 944188
rect 668252 943800 668328 944188
rect 159178 69900 159254 70200
rect 159366 69900 159442 70200
rect 161194 70153 161270 70200
rect 161194 70101 161206 70153
rect 161258 70101 161270 70153
rect 161194 69814 161270 70101
rect 162066 70055 162142 70200
rect 162066 70003 162079 70055
rect 162131 70003 162142 70055
rect 162066 69813 162142 70003
rect 174172 69813 174248 70200
rect 215672 70055 215748 70200
rect 215672 70003 215683 70055
rect 215735 70003 215748 70055
rect 215672 69813 215748 70003
rect 216193 70055 216269 70200
rect 216193 70003 216205 70055
rect 216257 70003 216269 70055
rect 216193 69813 216269 70003
rect 216422 70055 216498 70200
rect 216422 70003 216433 70055
rect 216485 70003 216498 70055
rect 216422 69813 216498 70003
rect 216564 70055 216640 70200
rect 216564 70003 216575 70055
rect 216627 70003 216640 70055
rect 216564 69813 216640 70003
rect 216706 69813 216782 70200
rect 217066 70055 217142 70200
rect 217066 70003 217077 70055
rect 217129 70003 217142 70055
rect 217066 69813 217142 70003
rect 217277 70055 217353 70200
rect 217277 70003 217289 70055
rect 217341 70003 217353 70055
rect 217277 69813 217353 70003
rect 228734 70055 228810 70200
rect 228734 70003 228746 70055
rect 228798 70003 228810 70055
rect 228734 69813 228810 70003
rect 228880 70055 228956 70200
rect 228880 70003 228891 70055
rect 228943 70003 228956 70055
rect 228880 69813 228956 70003
rect 229026 70055 229102 70200
rect 229026 70003 229037 70055
rect 229089 70003 229102 70055
rect 229026 69813 229102 70003
rect 229172 69813 229248 70200
rect 230558 69900 230634 70200
rect 230746 69900 230822 70200
rect 325672 69813 325748 70200
rect 326193 69813 326269 70200
rect 326422 69813 326498 70200
rect 326564 69813 326640 70200
rect 326706 69813 326782 70200
rect 327066 69813 327142 70200
rect 327277 69813 327353 70200
rect 338734 69813 338810 70200
rect 338880 69813 338956 70200
rect 339026 69813 339102 70200
rect 339172 69813 339248 70200
rect 340558 69900 340634 70200
rect 340746 69900 340822 70200
rect 380672 69813 380748 70200
rect 381193 69813 381269 70200
rect 381422 69813 381498 70200
rect 381564 69813 381640 70200
rect 381706 69813 381782 70200
rect 382066 69813 382142 70200
rect 382277 69813 382353 70200
rect 393734 69813 393810 70200
rect 393880 69813 393956 70200
rect 394026 69813 394102 70200
rect 394172 69813 394248 70200
rect 395558 69900 395634 70200
rect 395746 69900 395822 70200
rect 435672 69813 435748 70200
rect 436193 69813 436269 70200
rect 436422 69813 436498 70200
rect 436564 69813 436640 70200
rect 436706 69813 436782 70200
rect 437066 69813 437142 70200
rect 437277 69813 437353 70200
rect 448734 69813 448810 70200
rect 448880 69813 448956 70200
rect 449026 69813 449102 70200
rect 449171 69924 449248 70200
rect 449172 69813 449248 69924
rect 450558 69900 450634 70200
rect 450746 69900 450822 70200
rect 490672 69813 490748 70200
rect 491193 69813 491269 70200
rect 491422 69813 491498 70200
rect 491564 69813 491640 70200
rect 491706 69813 491782 70200
rect 492066 69813 492142 70200
rect 492277 69813 492353 70200
rect 503734 69813 503810 70200
rect 503880 69813 503956 70200
rect 504026 69813 504102 70200
rect 504172 69813 504248 70200
rect 505558 69900 505634 70200
rect 505746 69900 505822 70200
rect 507707 69900 507783 70200
rect 508290 69900 508366 70200
rect 509707 69900 509783 70200
rect 510290 69900 510366 70200
rect 511707 69900 511783 70200
rect 512290 69900 512366 70200
rect 513707 69900 513783 70200
rect 514290 69900 514366 70200
rect 515707 69900 515783 70200
rect 516290 69900 516366 70200
rect 517707 69900 517783 70200
rect 518290 69900 518366 70200
rect 519707 69900 519783 70200
rect 520290 69900 520366 70200
rect 521707 69900 521783 70200
rect 522290 69900 522366 70200
rect 523707 69900 523783 70200
rect 524290 69900 524366 70200
rect 525707 69900 525783 70200
rect 526290 69900 526366 70200
rect 527707 69900 527783 70200
rect 528290 69900 528366 70200
rect 529707 69900 529783 70200
rect 530290 69900 530366 70200
rect 531707 69900 531783 70200
rect 532290 69900 532366 70200
rect 533707 69900 533783 70200
rect 534290 69900 534366 70200
rect 535707 69900 535783 70200
rect 536290 69900 536366 70200
rect 537707 69900 537783 70200
rect 538290 69900 538366 70200
rect 507707 69848 507765 69900
rect 507707 69813 507763 69848
rect 508290 69813 508346 69900
rect 509707 69813 509763 69900
rect 510290 69813 510346 69900
rect 511707 69813 511763 69900
rect 512290 69813 512346 69900
rect 513707 69813 513763 69900
rect 514290 69813 514346 69900
rect 515707 69813 515763 69900
rect 516290 69813 516346 69900
rect 517707 69813 517763 69900
rect 518290 69813 518346 69900
rect 519707 69813 519763 69900
rect 520290 69813 520346 69900
rect 521707 69813 521763 69900
rect 522290 69813 522346 69900
rect 523707 69813 523763 69900
rect 524290 69813 524346 69900
rect 525707 69813 525763 69900
rect 526290 69813 526346 69900
rect 527707 69813 527763 69900
rect 528290 69813 528346 69900
rect 529707 69813 529763 69900
rect 530290 69813 530346 69900
rect 531707 69813 531763 69900
rect 532290 69813 532346 69900
rect 533707 69813 533763 69900
rect 534290 69813 534346 69900
rect 535707 69813 535763 69900
rect 536290 69813 536346 69900
rect 537707 69813 537763 69900
rect 538290 69813 538346 69900
rect 545672 69813 545748 70200
rect 546193 69813 546269 70200
rect 546422 69813 546498 70200
rect 546564 69813 546640 70200
rect 546706 69813 546782 70200
rect 547066 69813 547142 70200
rect 547277 69813 547353 70200
rect 558734 69813 558810 70200
rect 558880 69813 558956 70200
rect 559026 69813 559102 70200
rect 559172 69813 559248 70200
rect 560558 69900 560634 70200
rect 560746 69900 560822 70200
rect 590707 69900 590783 70200
rect 591290 69900 591366 70200
rect 593218 69900 593294 70200
rect 590707 69813 590763 69900
rect 591290 69813 591346 69900
rect 593218 69813 593274 69900
<< metal3 >>
rect 705729 921746 706029 921822
rect 705729 921558 706029 921634
rect 705729 920172 706005 920248
rect 705729 920026 706005 920102
rect 705729 919880 706005 919956
rect 705729 919734 706005 919810
rect 69995 919252 70271 919328
rect 69995 918731 70271 918807
rect 69995 918502 70271 918578
rect 69995 918360 70271 918436
rect 69995 918218 70271 918294
rect 69995 917858 70271 917934
rect 69995 917647 70271 917723
rect 705729 908277 706005 908353
rect 705729 908066 706005 908142
rect 705729 907706 706005 907782
rect 705729 907564 706005 907640
rect 705729 907422 706005 907498
rect 705729 907193 706005 907269
rect 705729 906672 706005 906748
rect 69995 906190 70271 906266
rect 69995 906044 70271 906120
rect 69995 905898 70271 905974
rect 69995 905752 70271 905828
rect 69971 904366 70271 904442
rect 69971 904178 70271 904254
rect 705729 835746 706029 835822
rect 705729 835558 706029 835634
rect 705729 834172 706005 834248
rect 705729 834026 706005 834102
rect 705729 833880 706005 833956
rect 705729 833734 706005 833810
rect 705729 822277 706005 822353
rect 705729 822066 706005 822142
rect 705729 821706 706005 821782
rect 705729 821564 706005 821640
rect 705729 821422 706005 821498
rect 705729 821193 706005 821269
rect 705729 820672 706005 820748
rect 69995 755252 70271 755328
rect 69995 754731 70271 754807
rect 69995 754502 70271 754578
rect 69995 754360 70271 754436
rect 69995 754218 70271 754294
rect 69995 753858 70271 753934
rect 69995 753647 70271 753723
rect 705729 749746 706029 749822
rect 705729 749558 706029 749634
rect 705729 748172 706005 748248
rect 705729 748026 706005 748102
rect 705729 747880 706005 747956
rect 705729 747734 706005 747810
rect 69995 742190 70271 742266
rect 69995 742044 70271 742120
rect 69995 741898 70271 741974
rect 69995 741752 70271 741828
rect 69971 740366 70271 740442
rect 69971 740178 70271 740254
rect 705729 736277 706005 736353
rect 705729 736066 706005 736142
rect 705729 735706 706005 735782
rect 705729 735564 706005 735640
rect 705729 735422 706005 735498
rect 705729 735193 706005 735269
rect 705729 734672 706005 734748
rect 69995 714252 70271 714328
rect 69995 713731 70271 713807
rect 69995 713502 70271 713578
rect 69995 713360 70271 713436
rect 69995 713218 70271 713294
rect 69995 712858 70271 712934
rect 69995 712647 70271 712723
rect 705729 706746 706029 706822
rect 705729 706558 706029 706634
rect 705729 705172 706005 705248
rect 705729 705026 706005 705102
rect 705729 704880 706005 704956
rect 705729 704734 706005 704810
rect 69995 701190 70271 701266
rect 69995 701044 70271 701120
rect 69995 700898 70271 700974
rect 69995 700752 70271 700828
rect 69971 699366 70271 699442
rect 69971 699178 70271 699254
rect 705729 693277 706005 693353
rect 705729 693066 706005 693142
rect 705729 692706 706005 692782
rect 705729 692564 706005 692640
rect 705729 692422 706005 692498
rect 705729 692193 706005 692269
rect 705729 691672 706005 691748
rect 69995 673252 70271 673328
rect 69995 672731 70271 672807
rect 69995 672502 70271 672578
rect 69995 672360 70271 672436
rect 69995 672218 70271 672294
rect 69995 671858 70271 671934
rect 69995 671647 70271 671723
rect 705729 663746 706029 663822
rect 705729 663558 706029 663634
rect 705729 662172 706005 662248
rect 705729 662026 706005 662102
rect 705729 661880 706005 661956
rect 705729 661734 706005 661810
rect 69995 660190 70271 660266
rect 69995 660044 70271 660120
rect 69995 659898 70271 659974
rect 69995 659752 70271 659828
rect 69971 658366 70271 658442
rect 69971 658178 70271 658254
rect 705729 650277 706005 650353
rect 705729 650066 706005 650142
rect 705729 649706 706005 649782
rect 705729 649564 706005 649640
rect 705729 649422 706005 649498
rect 705729 649193 706005 649269
rect 705729 648672 706005 648748
rect 69995 632252 70271 632328
rect 69995 631731 70271 631807
rect 69995 631502 70271 631578
rect 69995 631360 70271 631436
rect 69995 631218 70271 631294
rect 69995 630858 70271 630934
rect 69995 630647 70271 630723
rect 705729 620746 706029 620822
rect 705729 620558 706029 620634
rect 69995 619190 70271 619266
rect 705729 619172 706005 619248
rect 69995 619044 70271 619120
rect 705729 619026 706005 619102
rect 69995 618898 70271 618974
rect 705729 618880 706005 618956
rect 69995 618752 70271 618828
rect 705729 618734 706005 618810
rect 69971 617366 70271 617442
rect 69971 617178 70271 617254
rect 705729 607277 706005 607353
rect 705729 607066 706005 607142
rect 705729 606706 706005 606782
rect 705729 606564 706005 606640
rect 705729 606422 706005 606498
rect 705729 606193 706005 606269
rect 705729 605672 706005 605748
rect 69995 591252 70271 591328
rect 69995 590731 70271 590807
rect 69995 590502 70271 590578
rect 69995 590360 70271 590436
rect 69995 590218 70271 590294
rect 69995 589858 70271 589934
rect 69995 589647 70271 589723
rect 69995 578190 70271 578266
rect 69995 578044 70271 578120
rect 69995 577898 70271 577974
rect 69995 577752 70271 577828
rect 705729 577746 706029 577822
rect 705729 577558 706029 577634
rect 69971 576366 70271 576442
rect 69971 576178 70271 576254
rect 705729 576172 706005 576248
rect 705729 576026 706005 576102
rect 705729 575880 706005 575956
rect 705729 575734 706005 575810
rect 705729 564277 706005 564353
rect 705729 564066 706005 564142
rect 705729 563706 706005 563782
rect 705729 563564 706005 563640
rect 705729 563422 706005 563498
rect 705729 563193 706005 563269
rect 705729 562672 706005 562748
rect 69995 550252 70271 550328
rect 69995 549731 70271 549807
rect 69995 549502 70271 549578
rect 69995 549360 70271 549436
rect 69995 549218 70271 549294
rect 69995 548858 70271 548934
rect 69995 548647 70271 548723
rect 69995 537190 70271 537266
rect 69995 537044 70271 537120
rect 69995 536898 70271 536974
rect 69995 536752 70271 536828
rect 69971 535366 70271 535442
rect 69971 535178 70271 535254
rect 705729 534746 706029 534822
rect 705729 534558 706029 534634
rect 705729 533172 706005 533248
rect 705729 533026 706005 533102
rect 705729 532880 706005 532956
rect 705729 532734 706005 532810
rect 705729 521277 706005 521353
rect 705729 521066 706005 521142
rect 705729 520706 706005 520782
rect 705729 520564 706005 520640
rect 705729 520422 706005 520498
rect 705729 520193 706005 520269
rect 705729 519672 706005 519748
rect 69995 509252 70271 509328
rect 69995 508731 70271 508807
rect 69995 508502 70271 508578
rect 69995 508360 70271 508436
rect 69995 508218 70271 508294
rect 69995 507858 70271 507934
rect 69995 507647 70271 507723
rect 69995 496190 70271 496266
rect 69995 496044 70271 496120
rect 69995 495898 70271 495974
rect 69995 495752 70271 495828
rect 69971 494366 70271 494442
rect 69971 494178 70271 494254
rect 69995 386252 70271 386328
rect 69995 385731 70271 385807
rect 69995 385502 70271 385578
rect 69995 385360 70271 385436
rect 69995 385218 70271 385294
rect 69995 384858 70271 384934
rect 69995 384647 70271 384723
rect 69995 373190 70271 373266
rect 69995 373044 70271 373120
rect 69995 372898 70271 372974
rect 69995 372752 70271 372828
rect 69971 371366 70271 371442
rect 69971 371178 70271 371254
rect 705729 362746 706029 362822
rect 705729 362558 706029 362634
rect 705729 361172 706005 361248
rect 705729 361026 706005 361102
rect 705729 360880 706005 360956
rect 705729 360734 706005 360810
rect 705729 349277 706005 349353
rect 705729 349066 706005 349142
rect 705729 348706 706005 348782
rect 705729 348564 706005 348640
rect 705729 348422 706005 348498
rect 705729 348193 706005 348269
rect 705729 347672 706005 347748
rect 69995 345252 70271 345328
rect 69995 344731 70271 344807
rect 69995 344502 70271 344578
rect 69995 344360 70271 344436
rect 69995 344218 70271 344294
rect 69995 343858 70271 343934
rect 69995 343647 70271 343723
rect 69995 332190 70271 332266
rect 69995 332044 70271 332120
rect 69995 331898 70271 331974
rect 69995 331752 70271 331828
rect 69971 330366 70271 330442
rect 69971 330178 70271 330254
rect 705729 319746 706029 319822
rect 705729 319558 706029 319634
rect 705729 318172 706005 318248
rect 705729 318026 706005 318102
rect 705729 317880 706005 317956
rect 705729 317734 706005 317810
rect 705729 306277 706005 306353
rect 705729 306066 706005 306142
rect 705729 305706 706005 305782
rect 705729 305564 706005 305640
rect 705729 305422 706005 305498
rect 705729 305193 706005 305269
rect 705729 304672 706005 304748
rect 69995 304252 70271 304328
rect 69995 303731 70271 303807
rect 69995 303502 70271 303578
rect 69995 303360 70271 303436
rect 69995 303218 70271 303294
rect 69995 302858 70271 302934
rect 69995 302647 70271 302723
rect 69995 291190 70271 291266
rect 69995 291044 70271 291120
rect 69995 290898 70271 290974
rect 69995 290752 70271 290828
rect 69971 289366 70271 289442
rect 69971 289178 70271 289254
rect 705729 276746 706029 276822
rect 705729 276558 706029 276634
rect 705729 275172 706005 275248
rect 705729 275026 706005 275102
rect 705729 274880 706005 274956
rect 705729 274734 706005 274810
rect 69995 263252 70271 263328
rect 705729 263277 706005 263353
rect 705729 263066 706005 263142
rect 69995 262731 70271 262807
rect 705729 262706 706005 262782
rect 69995 262502 70271 262578
rect 705729 262564 706005 262640
rect 69995 262360 70271 262436
rect 705729 262422 706005 262498
rect 69995 262218 70271 262294
rect 705729 262193 706005 262269
rect 69995 261858 70271 261934
rect 69995 261647 70271 261723
rect 705729 261672 706005 261748
rect 69995 250190 70271 250266
rect 69995 250044 70271 250120
rect 69995 249898 70271 249974
rect 69995 249752 70271 249828
rect 69972 248366 70271 248442
rect 69972 248178 70271 248254
rect 705729 233746 706029 233822
rect 705729 233558 706029 233634
rect 705729 232172 706005 232248
rect 705729 232026 706005 232102
rect 705729 231880 706005 231956
rect 705729 231734 706005 231810
rect 69995 222252 70271 222328
rect 69995 221731 70271 221807
rect 69995 221502 70271 221578
rect 69995 221360 70271 221436
rect 69995 221218 70271 221294
rect 69995 220858 70271 220934
rect 69995 220647 70271 220723
rect 705729 220277 706005 220353
rect 705729 220066 706005 220142
rect 705729 219706 706005 219782
rect 705729 219564 706005 219640
rect 705729 219422 706005 219498
rect 705729 219193 706005 219269
rect 705729 218672 706005 218748
rect 69995 209190 70271 209266
rect 69995 209044 70271 209120
rect 69995 208898 70271 208974
rect 69995 208752 70271 208828
rect 69971 207366 70271 207442
rect 69971 207178 70271 207254
rect 705729 190746 706029 190822
rect 705729 190558 706029 190634
rect 705729 189172 706005 189248
rect 705729 189026 706005 189102
rect 705729 188880 706005 188956
rect 705729 188734 706005 188810
rect 69995 181252 70271 181328
rect 69995 180731 70271 180807
rect 69995 180502 70271 180578
rect 69995 180360 70271 180436
rect 69995 180218 70271 180294
rect 69995 179858 70271 179934
rect 69995 179647 70271 179723
rect 705729 177277 706005 177353
rect 705729 177066 706005 177142
rect 705729 176706 706005 176782
rect 705729 176564 706005 176640
rect 705729 176422 706005 176498
rect 705729 176193 706005 176269
rect 705729 175672 706005 175748
rect 69995 168190 70271 168266
rect 69995 168044 70271 168120
rect 69995 167898 70271 167974
rect 69995 167752 70271 167828
rect 69971 166366 70271 166442
rect 69971 166178 70271 166254
rect 705729 147746 706029 147822
rect 705729 147558 706029 147634
rect 705729 146172 706119 146248
rect 705729 146026 706119 146102
rect 705729 145880 706119 145956
rect 705729 145734 706119 145810
rect 705729 134277 706128 134353
rect 705729 134066 706128 134142
rect 705729 133706 706107 133782
rect 705729 133564 706128 133640
rect 705729 133422 706128 133498
rect 705729 133193 706128 133269
rect 705729 132672 706128 132748
rect 705729 104746 706029 104822
rect 705729 104558 706029 104634
rect 705729 103172 706005 103248
rect 705729 103026 706005 103102
rect 705729 102880 706005 102956
rect 705729 102734 706005 102810
rect 705729 91277 706005 91353
rect 705729 91066 706005 91142
rect 705729 90706 706005 90782
rect 705729 90564 706005 90640
rect 705729 90422 706005 90498
rect 705729 90193 706005 90269
rect 705729 89672 706005 89748
<< metal4 >>
rect 379272 943800 381172 944000
rect 381752 943800 383802 944000
rect 384122 943800 386172 944000
rect 386828 943800 388878 944000
rect 389198 943800 391248 944000
rect 391828 943800 393728 944000
rect 599272 943800 601172 944000
rect 601752 943800 603802 944000
rect 604122 943800 606172 944000
rect 606828 943800 608878 944000
rect 609198 943800 611248 944000
rect 611828 943800 613728 944000
rect 105272 70000 107172 70200
rect 107752 70000 109802 70200
rect 110122 70000 112172 70200
rect 112828 70000 114878 70200
rect 115198 70000 117248 70200
rect 117828 70000 119728 70200
rect 270272 70000 272172 70200
rect 272752 70000 274802 70200
rect 275122 70000 277172 70200
rect 277828 70000 279878 70200
rect 280198 70000 282248 70200
rect 282828 70000 284728 70200
rect 600272 70000 602172 70200
rect 602752 70000 604802 70200
rect 605122 70000 607172 70200
rect 607828 70000 609878 70200
rect 610198 70000 612248 70200
rect 612828 70000 614728 70200
rect 655272 69999 657172 70199
rect 657752 69999 659802 70199
rect 660122 69999 662172 70199
rect 662828 69999 664878 70199
rect 665198 69999 667248 70199
rect 667828 69999 669728 70199
<< metal5 >>
rect 70000 876828 70270 878728
rect 70000 874198 70270 876248
rect 705730 875828 706000 877728
rect 70000 871828 70270 873878
rect 705728 873186 706002 875260
rect 70000 869122 70270 871172
rect 705730 870828 706000 872878
rect 70000 866752 70270 868802
rect 705728 868110 706002 870184
rect 70000 864272 70270 866172
rect 705730 865752 706000 867802
rect 705728 863260 706002 865184
rect 70000 835828 70270 837728
rect 70000 833198 70270 835248
rect 70000 830828 70270 832878
rect 70000 828122 70270 830172
rect 70000 825752 70270 827802
rect 70000 823272 70270 825172
rect 70000 794829 70270 796729
rect 70000 792199 70270 794249
rect 70000 789829 70270 791879
rect 705730 789828 706000 791728
rect 70000 787123 70270 789173
rect 705728 787186 706002 789260
rect 70000 784753 70270 786803
rect 705730 784828 706000 786878
rect 70000 782273 70270 784173
rect 705728 782110 706002 784184
rect 705730 779752 706000 781802
rect 705726 777248 706004 779196
rect 705730 488828 706000 490728
rect 705730 486198 706000 488248
rect 705730 483828 706000 485878
rect 705730 481122 706000 483172
rect 705730 478752 706000 480802
rect 705730 476272 706000 478172
rect 70000 466828 70270 468728
rect 70000 464198 70270 466248
rect 70000 461828 70270 463878
rect 70000 459122 70270 461172
rect 70000 456752 70270 458802
rect 70000 454272 70270 456172
rect 705730 445828 706000 447728
rect 705730 443198 706000 445248
rect 705730 440828 706000 442878
rect 705730 438122 706000 440172
rect 705730 435752 706000 437802
rect 705730 433272 706000 435172
rect 70000 425828 70270 427728
rect 69998 423186 70272 425260
rect 70000 420828 70270 422878
rect 70000 418122 70270 420172
rect 69998 415740 70272 417814
rect 70000 413272 70270 415172
rect 705730 402828 706000 404728
rect 705730 400198 706000 402248
rect 705730 397828 706000 399878
rect 705730 395122 706000 397172
rect 705730 392752 706000 394802
rect 705730 390272 706000 392172
rect 70000 138828 70270 140728
rect 69998 136186 70272 138260
rect 70000 133828 70270 135878
rect 70000 131122 70270 133172
rect 69998 128740 70272 130814
rect 70000 126272 70270 128172
rect 70000 97828 70270 99728
rect 69998 95186 70272 97260
rect 70000 92828 70270 94878
rect 70000 90122 70270 92172
rect 69998 87740 70272 89814
rect 70000 85272 70270 87172
<< comment >>
rect 69593 944007 706407 944407
rect 69593 69993 69993 944007
rect 70013 943983 705987 943987
rect 70013 70017 70017 943983
rect 705983 70017 705987 943983
rect 70013 70013 705987 70017
rect 706007 69993 706407 944007
rect 69593 69593 706407 69993
use horz_connects_gpio_disabled  horz_connects_gpio_disabled_1
timestamp 1764975181
transform 1 0 215490 0 1 69968
box 0 0 15507 232
use horz_connects_gpio_disabled  horz_connects_gpio_disabled_2
timestamp 1764975181
transform 1 0 325490 0 1 69968
box 0 0 15507 232
use horz_connects_gpio_disabled  horz_connects_gpio_disabled_3
timestamp 1764975181
transform 1 0 380490 0 1 69968
box 0 0 15507 232
use horz_connects_gpio_disabled  horz_connects_gpio_disabled_4
timestamp 1764975181
transform 1 0 435490 0 1 69968
box 0 0 15507 232
use horz_connects_gpio_disabled  horz_connects_gpio_disabled_5
timestamp 1764975181
transform 1 0 490490 0 1 69968
box 0 0 15507 232
use horz_connects_gpio_disabled  horz_connects_gpio_disabled_6
timestamp 1764975181
transform 1 0 545490 0 1 69968
box 0 0 15507 232
use horz_connects_gpio_disabled  horz_connects_gpio_disabled_7
timestamp 1764975181
transform -1 0 668510 0 -1 944032
box 0 0 15507 232
use horz_connects_gpio_disabled  horz_connects_gpio_disabled_8
timestamp 1764975181
transform -1 0 558510 0 -1 944032
box 0 0 15507 232
use horz_connects_gpio_disabled  horz_connects_gpio_disabled_9
timestamp 1764975181
transform -1 0 503510 0 -1 944032
box 0 0 15507 232
use horz_connects_gpio_disabled  horz_connects_gpio_disabled_10
timestamp 1764975181
transform -1 0 448510 0 -1 944032
box 0 0 15507 232
use horz_connects_gpio_disabled  horz_connects_gpio_disabled_11
timestamp 1764975181
transform -1 0 338510 0 -1 944032
box 0 0 15507 232
use horz_connects_gpio_disabled  horz_connects_gpio_disabled_12
timestamp 1764975181
transform -1 0 283510 0 -1 944032
box 0 0 15507 232
use horz_connects_gpio_disabled  horz_connects_gpio_disabled_13
timestamp 1764975181
transform -1 0 228510 0 -1 944032
box 0 0 15507 232
use horz_connects_gpio_disabled  horz_connects_gpio_disabled_14
timestamp 1764975181
transform -1 0 173510 0 -1 944032
box 0 0 15507 232
use horz_connects_gpio_disabled  horz_connects_gpio_disabled_15
timestamp 1764975181
transform -1 0 118510 0 -1 944032
box 0 0 15507 232
use horz_connects_resetb_pullup  horz_connects_resetb_pullup_0
timestamp 1764982896
transform 1 0 159058 0 1 69968
box -75 0 3129 232
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_0
timestamp 1764982451
transform 1 0 69968 0 1 166058
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_1
timestamp 1764982451
transform 1 0 69968 0 1 207058
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_2
timestamp 1764982451
transform 1 0 69968 0 1 289058
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_3
timestamp 1764982451
transform 1 0 69968 0 1 330058
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_4
timestamp 1764982451
transform 1 0 69968 0 1 371058
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_5
timestamp 1764982451
transform 1 0 69968 0 1 494058
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_6
timestamp 1764982451
transform 1 0 69968 0 1 535058
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_7
timestamp 1764982451
transform 1 0 69968 0 1 576058
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_8
timestamp 1764982451
transform 1 0 69968 0 1 617058
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_9
timestamp 1764982451
transform 1 0 69968 0 1 658058
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_10
timestamp 1764982451
transform 1 0 69968 0 1 699058
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_11
timestamp 1764982451
transform 1 0 69968 0 1 740058
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_12
timestamp 1764982451
transform 1 0 69968 0 1 904058
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_13
timestamp 1764982451
transform -1 0 706032 0 -1 104942
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_14
timestamp 1764982451
transform -1 0 706032 0 -1 147942
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_15
timestamp 1764982451
transform -1 0 706032 0 -1 190942
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_16
timestamp 1764982451
transform -1 0 706032 0 -1 233942
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_17
timestamp 1764982451
transform -1 0 706032 0 -1 276942
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_18
timestamp 1764982451
transform -1 0 706032 0 -1 319942
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_19
timestamp 1764982451
transform -1 0 706032 0 -1 362942
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_20
timestamp 1764982451
transform -1 0 706032 0 -1 534942
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_21
timestamp 1764982451
transform -1 0 706032 0 -1 577942
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_22
timestamp 1764982451
transform -1 0 706032 0 -1 620942
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_23
timestamp 1764982451
transform -1 0 706032 0 -1 663942
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_24
timestamp 1764982451
transform -1 0 706032 0 -1 706942
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_25
timestamp 1764982451
transform -1 0 706032 0 -1 749942
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_26
timestamp 1764982451
transform -1 0 706032 0 -1 835942
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_27
timestamp 1764982451
transform -1 0 706032 0 -1 921942
box 0 -6 303 15452
use vert_connects_gpio_disabled  vert_connects_gpio_disabled_28
timestamp 1764982451
transform 1 0 69968 0 1 248058
box 0 -6 303 15452
<< labels >>
flabel metal2 505558 69900 505634 70200 0 FreeSans 480 90 0 0 gpio_loopback_one[42]
port 582 nsew
flabel metal2 505746 69900 505822 70200 0 FreeSans 480 90 0 0 gpio_loopback_zero[42]
port 581 nsew
flabel metal2 395558 69900 395634 70200 0 FreeSans 480 90 0 0 gpio_loopback_one[40]
port 578 nsew
flabel metal2 395746 69900 395822 70200 0 FreeSans 480 90 0 0 gpio_loopback_zero[40]
port 577 nsew
flabel metal2 230558 69900 230634 70200 0 FreeSans 480 90 0 0 gpio_loopback_one[38]
port 573 nsew
flabel metal2 230746 69900 230822 70200 0 FreeSans 480 90 0 0 gpio_loopback_zero[38]
port 572 nsew
flabel metal2 103178 943800 103254 944100 0 FreeSans 480 90 0 0 gpio_loopback_zero[23]
port 543 nsew
flabel metal2 103366 943800 103442 944100 0 FreeSans 480 90 0 0 gpio_loopback_one[23]
port 542 nsew
flabel metal2 213178 943800 213254 944100 0 FreeSans 480 90 0 0 gpio_loopback_zero[21]
port 539 nsew
flabel metal2 213366 943800 213442 944100 0 FreeSans 480 90 0 0 gpio_loopback_one[21]
port 538 nsew
flabel metal2 323178 943800 323254 944100 0 FreeSans 480 90 0 0 gpio_loopback_zero[19]
port 535 nsew
flabel metal2 323366 943800 323442 944100 0 FreeSans 480 90 0 0 gpio_loopback_one[19]
port 534 nsew
flabel metal2 488178 943800 488254 944100 0 FreeSans 480 90 0 0 gpio_loopback_zero[17]
port 531 nsew
flabel metal2 488366 943800 488442 944100 0 FreeSans 480 90 0 0 gpio_loopback_one[17]
port 530 nsew
flabel metal2 229026 69924 229102 70200 0 FreeSans 480 90 0 0 gpio_oe[38]
port 24 nsew
flabel metal2 228880 69924 228956 70200 0 FreeSans 480 90 0 0 gpio_out[38]
port 23 nsew
flabel metal2 228734 69924 228810 70200 0 FreeSans 480 90 0 0 gpio_slew[38]
port 28 nsew
flabel metal2 217277 69924 217353 70200 0 FreeSans 480 90 0 0 gpio_ie[38]
port 22 nsew
flabel metal2 217066 69924 217142 70200 0 FreeSans 480 90 0 0 gpio_pulldown[38]
port 25 nsew
flabel metal2 216706 69923 216782 70199 0 FreeSans 480 90 0 0 gpio_ana[38]
port 490 nsew
flabel metal2 216193 69924 216269 70200 0 FreeSans 480 90 0 0 gpio_pullup[38]
port 26 nsew
flabel metal2 216564 69923 216640 70199 0 FreeSans 480 90 0 0 gpio_drive1[38]
port 20 nsew
flabel metal2 216422 69924 216498 70200 0 FreeSans 480 90 0 0 gpio_drive0[38]
port 19 nsew
flabel metal2 215672 69924 215748 70200 0 FreeSans 480 90 0 0 gpio_schmitt[38]
port 27 nsew
flabel metal2 229172 69924 229248 70200 0 FreeSans 480 90 0 0 gpio_in[38]
port 1 nsew
flabel metal2 490672 69924 490748 70200 0 FreeSans 480 90 0 0 gpio_schmitt[42]
port 29 nsew
flabel metal2 491193 69924 491269 70200 0 FreeSans 480 90 0 0 gpio_pullup[42]
port 30 nsew
flabel metal2 491422 69924 491498 70200 0 FreeSans 480 90 0 0 gpio_drive0[42]
port 31 nsew
flabel metal2 491564 69923 491640 70199 0 FreeSans 480 90 0 0 gpio_drive1[42]
port 32 nsew
flabel metal2 491706 69923 491782 70199 0 FreeSans 480 90 0 0 gpio_ana[42]
port 494 nsew
flabel metal2 492066 69924 492142 70200 0 FreeSans 480 90 0 0 gpio_pulldown[42]
port 33 nsew
flabel metal2 503734 69924 503810 70200 0 FreeSans 480 90 0 0 gpio_slew[42]
port 34 nsew
flabel metal2 435672 69924 435748 70200 0 FreeSans 480 90 0 0 gpio_schmitt[41]
port 35 nsew
flabel metal2 436193 69924 436269 70200 0 FreeSans 480 90 0 0 gpio_pullup[41]
port 36 nsew
flabel metal2 436422 69924 436498 70200 0 FreeSans 480 90 0 0 gpio_drive0[41]
port 37 nsew
flabel metal2 436564 69923 436640 70199 0 FreeSans 480 90 0 0 gpio_drive1[41]
port 38 nsew
flabel metal2 436706 69923 436782 70199 0 FreeSans 480 90 0 0 gpio_ana[41]
port 493 nsew
flabel metal2 437066 69924 437142 70200 0 FreeSans 480 90 0 0 gpio_pulldown[41]
port 39 nsew
flabel metal2 448734 69924 448810 70200 0 FreeSans 480 90 0 0 gpio_slew[41]
port 40 nsew
flabel metal2 380672 69924 380748 70200 0 FreeSans 480 90 0 0 gpio_schmitt[40]
port 41 nsew
flabel metal2 381193 69924 381269 70200 0 FreeSans 480 90 0 0 gpio_pullup[40]
port 42 nsew
flabel metal2 381422 69924 381498 70200 0 FreeSans 480 90 0 0 gpio_drive0[40]
port 43 nsew
flabel metal2 381564 69923 381640 70199 0 FreeSans 480 90 0 0 gpio_drive1[40]
port 44 nsew
flabel metal2 381706 69923 381782 70199 0 FreeSans 480 90 0 0 gpio_ana[40]
port 492 nsew
flabel metal2 382066 69924 382142 70200 0 FreeSans 480 90 0 0 gpio_pulldown[40]
port 45 nsew
flabel metal2 382277 69924 382353 70200 0 FreeSans 480 90 0 0 gpio_ie[40]
port 46 nsew
flabel metal2 393734 69924 393810 70200 0 FreeSans 480 90 0 0 gpio_slew[40]
port 47 nsew
flabel metal2 393880 69924 393956 70200 0 FreeSans 480 90 0 0 gpio_out[40]
port 48 nsew
flabel metal2 325672 69924 325748 70200 0 FreeSans 480 90 0 0 gpio_schmitt[39]
port 49 nsew
flabel metal2 326193 69924 326269 70200 0 FreeSans 480 90 0 0 gpio_pullup[39]
port 50 nsew
flabel metal2 326422 69924 326498 70200 0 FreeSans 480 90 0 0 gpio_drive0[39]
port 51 nsew
flabel metal2 326564 69923 326640 70199 0 FreeSans 480 90 0 0 gpio_drive1[39]
port 52 nsew
flabel metal2 326706 69923 326782 70199 0 FreeSans 480 90 0 0 gpio_ana[39]
port 491 nsew
flabel metal2 327066 69924 327142 70200 0 FreeSans 480 90 0 0 gpio_pulldown[39]
port 53 nsew
flabel metal2 327277 69924 327353 70200 0 FreeSans 480 90 0 0 gpio_ie[39]
port 54 nsew
flabel metal2 338734 69924 338810 70200 0 FreeSans 480 90 0 0 gpio_slew[39]
port 55 nsew
flabel metal2 338880 69924 338956 70200 0 FreeSans 480 90 0 0 gpio_out[39]
port 56 nsew
flabel metal2 339026 69924 339102 70200 0 FreeSans 480 90 0 0 gpio_oe[39]
port 7 nsew
flabel metal2 339172 69924 339248 70200 0 FreeSans 480 90 0 0 gpio_in[39]
port 6 nsew
flabel metal2 394026 69924 394102 70200 0 FreeSans 480 90 0 0 gpio_oe[40]
port 4 nsew
flabel metal2 394172 69924 394248 70200 0 FreeSans 480 90 0 0 gpio_in[40]
port 3 nsew
flabel metal2 546706 69923 546782 70199 0 FreeSans 480 90 0 0 gpio_ana[43]
port 495 nsew
flabel metal2 117218 943800 117294 944076 0 FreeSans 480 270 0 0 gpio_ana[23]
port 475 nsew
flabel metal2 172218 943800 172294 944076 0 FreeSans 480 270 0 0 gpio_ana[22]
port 474 nsew
flabel metal2 227218 943800 227294 944076 0 FreeSans 480 270 0 0 gpio_ana[21]
port 473 nsew
flabel metal2 282218 943800 282294 944076 0 FreeSans 480 270 0 0 gpio_ana[20]
port 472 nsew
flabel metal2 337218 943800 337294 944076 0 FreeSans 480 270 0 0 gpio_ana[19]
port 471 nsew
flabel metal2 447218 943800 447294 944076 0 FreeSans 480 270 0 0 gpio_ana[18]
port 470 nsew
flabel metal2 502218 943800 502294 944076 0 FreeSans 480 270 0 0 gpio_ana[17]
port 469 nsew
flabel metal2 557218 943800 557294 944076 0 FreeSans 480 270 0 0 gpio_ana[16]
port 468 nsew
flabel metal2 667218 943800 667294 944076 0 FreeSans 480 270 0 0 gpio_ana[15]
port 467 nsew
flabel metal2 104752 943800 104828 944076 0 FreeSans 480 270 0 0 gpio_in[23]
port 157 nsew
flabel metal2 104898 943800 104974 944076 0 FreeSans 480 270 0 0 gpio_oe[23]
port 271 nsew
flabel metal2 105044 943800 105120 944076 0 FreeSans 480 270 0 0 gpio_out[23]
port 233 nsew
flabel metal2 105190 943800 105266 944076 0 FreeSans 480 270 0 0 gpio_slew[23]
port 423 nsew
flabel metal2 116647 943800 116723 944076 0 FreeSans 480 270 0 0 gpio_ie[23]
port 195 nsew
flabel metal2 116858 943800 116934 944076 0 FreeSans 480 270 0 0 gpio_pulldown[23]
port 309 nsew
flabel metal2 117360 943800 117436 944076 0 FreeSans 480 270 0 0 gpio_drive1[23]
port 108 nsew
flabel metal2 117502 943800 117578 944076 0 FreeSans 480 270 0 0 gpio_drive0[23]
port 107 nsew
flabel metal2 117731 943800 117807 944076 0 FreeSans 480 270 0 0 gpio_pullup[23]
port 347 nsew
flabel metal2 118252 943800 118328 944076 0 FreeSans 480 270 0 0 gpio_schmitt[23]
port 385 nsew
flabel metal2 159752 943800 159828 944076 0 FreeSans 480 270 0 0 gpio_in[22]
port 156 nsew
flabel metal2 159898 943800 159974 944076 0 FreeSans 480 270 0 0 gpio_oe[22]
port 270 nsew
flabel metal2 160044 943800 160120 944076 0 FreeSans 480 270 0 0 gpio_out[22]
port 232 nsew
flabel metal2 160190 943800 160266 944076 0 FreeSans 480 270 0 0 gpio_slew[22]
port 422 nsew
flabel metal2 171647 943800 171723 944076 0 FreeSans 480 270 0 0 gpio_ie[22]
port 194 nsew
flabel metal2 171858 943800 171934 944076 0 FreeSans 480 270 0 0 gpio_pulldown[22]
port 308 nsew
flabel metal2 172360 943800 172436 944076 0 FreeSans 480 270 0 0 gpio_drive1[22]
port 106 nsew
flabel metal2 172502 943800 172578 944076 0 FreeSans 480 270 0 0 gpio_drive0[22]
port 105 nsew
flabel metal2 172731 943800 172807 944076 0 FreeSans 480 270 0 0 gpio_pullup[22]
port 346 nsew
flabel metal2 173252 943800 173328 944076 0 FreeSans 480 270 0 0 gpio_schmitt[22]
port 384 nsew
flabel metal2 214752 943800 214828 944076 0 FreeSans 480 270 0 0 gpio_in[21]
port 155 nsew
flabel metal2 214898 943800 214974 944076 0 FreeSans 480 270 0 0 gpio_oe[21]
port 269 nsew
flabel metal2 215044 943800 215120 944076 0 FreeSans 480 270 0 0 gpio_out[21]
port 231 nsew
flabel metal2 215190 943800 215266 944076 0 FreeSans 480 270 0 0 gpio_slew[21]
port 421 nsew
flabel metal2 226647 943800 226723 944076 0 FreeSans 480 270 0 0 gpio_ie[21]
port 193 nsew
flabel metal2 226858 943800 226934 944076 0 FreeSans 480 270 0 0 gpio_pulldown[21]
port 307 nsew
flabel metal2 227360 943800 227436 944076 0 FreeSans 480 270 0 0 gpio_drive1[21]
port 104 nsew
flabel metal2 227502 943800 227578 944076 0 FreeSans 480 270 0 0 gpio_drive0[21]
port 103 nsew
flabel metal2 227731 943800 227807 944076 0 FreeSans 480 270 0 0 gpio_pullup[21]
port 345 nsew
flabel metal2 228252 943800 228328 944076 0 FreeSans 480 270 0 0 gpio_schmitt[21]
port 383 nsew
flabel metal2 269752 943800 269828 944076 0 FreeSans 480 270 0 0 gpio_in[20]
port 154 nsew
flabel metal2 269898 943800 269974 944076 0 FreeSans 480 270 0 0 gpio_oe[20]
port 268 nsew
flabel metal2 270044 943800 270120 944076 0 FreeSans 480 270 0 0 gpio_out[20]
port 230 nsew
flabel metal2 270190 943800 270266 944076 0 FreeSans 480 270 0 0 gpio_slew[20]
port 420 nsew
flabel metal2 281647 943800 281723 944076 0 FreeSans 480 270 0 0 gpio_ie[20]
port 192 nsew
flabel metal2 281858 943800 281934 944076 0 FreeSans 480 270 0 0 gpio_pulldown[20]
port 306 nsew
flabel metal2 282360 943800 282436 944076 0 FreeSans 480 270 0 0 gpio_drive1[20]
port 102 nsew
flabel metal2 282502 943800 282578 944076 0 FreeSans 480 270 0 0 gpio_drive0[20]
port 101 nsew
flabel metal2 282731 943800 282807 944076 0 FreeSans 480 270 0 0 gpio_pullup[20]
port 344 nsew
flabel metal2 283252 943800 283328 944076 0 FreeSans 480 270 0 0 gpio_schmitt[20]
port 382 nsew
flabel metal2 324752 943800 324828 944076 0 FreeSans 480 270 0 0 gpio_in[19]
port 152 nsew
flabel metal2 324898 943800 324974 944076 0 FreeSans 480 270 0 0 gpio_oe[19]
port 266 nsew
flabel metal2 325044 943800 325120 944076 0 FreeSans 480 270 0 0 gpio_out[19]
port 228 nsew
flabel metal2 325190 943800 325266 944076 0 FreeSans 480 270 0 0 gpio_slew[19]
port 418 nsew
flabel metal2 336647 943800 336723 944076 0 FreeSans 480 270 0 0 gpio_ie[19]
port 190 nsew
flabel metal2 336858 943800 336934 944076 0 FreeSans 480 270 0 0 gpio_pulldown[19]
port 304 nsew
flabel metal2 337360 943800 337436 944076 0 FreeSans 480 270 0 0 gpio_drive1[19]
port 99 nsew
flabel metal2 337502 943800 337578 944076 0 FreeSans 480 270 0 0 gpio_drive0[19]
port 98 nsew
flabel metal2 337731 943800 337807 944076 0 FreeSans 480 270 0 0 gpio_pullup[19]
port 342 nsew
flabel metal2 338252 943800 338328 944076 0 FreeSans 480 270 0 0 gpio_schmitt[19]
port 380 nsew
flabel metal2 434752 943800 434828 944076 0 FreeSans 480 270 0 0 gpio_in[18]
port 151 nsew
flabel metal2 434898 943800 434974 944076 0 FreeSans 480 270 0 0 gpio_oe[18]
port 265 nsew
flabel metal2 435044 943800 435120 944076 0 FreeSans 480 270 0 0 gpio_out[18]
port 227 nsew
flabel metal2 435190 943800 435266 944076 0 FreeSans 480 270 0 0 gpio_slew[18]
port 417 nsew
flabel metal2 446647 943800 446723 944076 0 FreeSans 480 270 0 0 gpio_ie[18]
port 189 nsew
flabel metal2 446858 943800 446934 944076 0 FreeSans 480 270 0 0 gpio_pulldown[18]
port 303 nsew
flabel metal2 447360 943800 447436 944076 0 FreeSans 480 270 0 0 gpio_drive1[18]
port 97 nsew
flabel metal2 447502 943800 447578 944076 0 FreeSans 480 270 0 0 gpio_drive0[18]
port 96 nsew
flabel metal2 447731 943800 447807 944076 0 FreeSans 480 270 0 0 gpio_pullup[18]
port 341 nsew
flabel metal2 448252 943800 448328 944076 0 FreeSans 480 270 0 0 gpio_schmitt[18]
port 379 nsew
flabel metal2 489752 943800 489828 944076 0 FreeSans 480 270 0 0 gpio_in[17]
port 150 nsew
flabel metal2 489898 943800 489974 944076 0 FreeSans 480 270 0 0 gpio_oe[17]
port 264 nsew
flabel metal2 490044 943800 490120 944076 0 FreeSans 480 270 0 0 gpio_out[17]
port 226 nsew
flabel metal2 490190 943800 490266 944076 0 FreeSans 480 270 0 0 gpio_slew[17]
port 416 nsew
flabel metal2 501647 943800 501723 944076 0 FreeSans 480 270 0 0 gpio_ie[17]
port 188 nsew
flabel metal2 501858 943800 501934 944076 0 FreeSans 480 270 0 0 gpio_pulldown[17]
port 302 nsew
flabel metal2 502360 943800 502436 944076 0 FreeSans 480 270 0 0 gpio_drive1[17]
port 95 nsew
flabel metal2 502502 943800 502578 944076 0 FreeSans 480 270 0 0 gpio_drive0[17]
port 94 nsew
flabel metal2 502731 943800 502807 944076 0 FreeSans 480 270 0 0 gpio_pullup[17]
port 340 nsew
flabel metal2 503252 943800 503328 944076 0 FreeSans 480 270 0 0 gpio_schmitt[17]
port 378 nsew
flabel metal2 544752 943800 544828 944076 0 FreeSans 480 270 0 0 gpio_in[16]
port 149 nsew
flabel metal2 544898 943800 544974 944076 0 FreeSans 480 270 0 0 gpio_oe[16]
port 263 nsew
flabel metal2 545044 943800 545120 944076 0 FreeSans 480 270 0 0 gpio_out[16]
port 225 nsew
flabel metal2 545190 943800 545266 944076 0 FreeSans 480 270 0 0 gpio_slew[16]
port 415 nsew
flabel metal2 556647 943800 556723 944076 0 FreeSans 480 270 0 0 gpio_ie[16]
port 187 nsew
flabel metal2 556858 943800 556934 944076 0 FreeSans 480 270 0 0 gpio_pulldown[16]
port 301 nsew
flabel metal2 557360 943800 557436 944076 0 FreeSans 480 270 0 0 gpio_drive1[16]
port 93 nsew
flabel metal2 557502 943800 557578 944076 0 FreeSans 480 270 0 0 gpio_drive0[16]
port 92 nsew
flabel metal2 557731 943800 557807 944076 0 FreeSans 480 270 0 0 gpio_pullup[16]
port 339 nsew
flabel metal2 558252 943800 558328 944076 0 FreeSans 480 270 0 0 gpio_schmitt[16]
port 377 nsew
flabel metal2 654752 943800 654828 944076 0 FreeSans 480 270 0 0 gpio_in[15]
port 148 nsew
flabel metal2 654898 943800 654974 944076 0 FreeSans 480 270 0 0 gpio_oe[15]
port 262 nsew
flabel metal2 655044 943800 655120 944076 0 FreeSans 480 270 0 0 gpio_out[15]
port 224 nsew
flabel metal2 655190 943800 655266 944076 0 FreeSans 480 270 0 0 gpio_slew[15]
port 414 nsew
flabel metal2 666647 943800 666723 944076 0 FreeSans 480 270 0 0 gpio_ie[15]
port 186 nsew
flabel metal2 666858 943800 666934 944076 0 FreeSans 480 270 0 0 gpio_pulldown[15]
port 300 nsew
flabel metal2 667360 943800 667436 944076 0 FreeSans 480 270 0 0 gpio_drive1[15]
port 91 nsew
flabel metal2 667502 943800 667578 944076 0 FreeSans 480 270 0 0 gpio_drive0[15]
port 90 nsew
flabel metal2 667731 943800 667807 944076 0 FreeSans 480 270 0 0 gpio_pullup[15]
port 338 nsew
flabel metal2 668252 943800 668328 944076 0 FreeSans 480 270 0 0 gpio_schmitt[15]
port 376 nsew
flabel metal2 559026 69924 559102 70200 0 FreeSans 480 90 0 0 gpio_oe[43]
port 65 nsew
flabel metal2 559172 69924 559248 70200 0 FreeSans 480 90 0 0 gpio_in[43]
port 21 nsew
flabel metal2 558880 69924 558956 70200 0 FreeSans 480 90 0 0 gpio_out[43]
port 57 nsew
flabel metal2 558734 69924 558810 70200 0 FreeSans 480 90 0 0 gpio_slew[43]
port 58 nsew
flabel metal2 547277 69924 547353 70200 0 FreeSans 480 90 0 0 gpio_ie[43]
port 59 nsew
flabel metal2 547066 69924 547142 70200 0 FreeSans 480 90 0 0 gpio_pulldown[43]
port 60 nsew
flabel metal2 546564 69923 546640 70199 0 FreeSans 480 90 0 0 gpio_drive1[43]
port 61 nsew
flabel metal2 546422 69924 546498 70200 0 FreeSans 480 90 0 0 gpio_drive0[43]
port 62 nsew
flabel metal2 546193 69924 546269 70200 0 FreeSans 480 90 0 0 gpio_pullup[43]
port 63 nsew
flabel metal2 545672 69924 545748 70200 0 FreeSans 480 90 0 0 gpio_schmitt[43]
port 64 nsew
flabel metal2 504172 69924 504248 70200 0 FreeSans 480 90 0 0 gpio_in[42]
port 14 nsew
flabel metal2 504026 69924 504102 70200 0 FreeSans 480 90 0 0 gpio_oe[42]
port 17 nsew
flabel metal2 503880 69924 503956 70200 0 FreeSans 480 90 0 0 gpio_out[42]
port 15 nsew
flabel metal2 492277 69924 492353 70200 0 FreeSans 480 90 0 0 gpio_ie[42]
port 16 nsew
flabel metal2 449171 69924 449247 70200 0 FreeSans 480 90 0 0 gpio_in[41]
port 9 nsew
flabel metal2 449026 69924 449102 70200 0 FreeSans 480 90 0 0 gpio_oe[41]
port 12 nsew
flabel metal2 448880 69924 448956 70200 0 FreeSans 480 90 0 0 gpio_out[41]
port 10 nsew
flabel metal2 437277 69924 437353 70200 0 FreeSans 480 90 0 0 gpio_ie[41]
port 11 nsew
flabel metal2 174172 69924 174248 70200 0 FreeSans 480 90 0 0 resetb_core
port 447 nsew
flabel metal3 705730 146172 706006 146248 0 FreeSans 480 0 0 0 gpio_in[1]
port 153 nsew
flabel metal3 705730 146026 706006 146102 0 FreeSans 480 0 0 0 gpio_oe[1]
port 267 nsew
flabel metal3 705730 145880 706006 145956 0 FreeSans 480 0 0 0 gpio_out[1]
port 229 nsew
flabel metal3 705730 145734 706006 145810 0 FreeSans 480 0 0 0 gpio_slew[1]
port 419 nsew
flabel metal3 705729 133706 706005 133782 0 FreeSans 480 0 0 0 gpio_ana[1]
port 453 nsew
flabel metal3 705729 133564 706005 133640 0 FreeSans 480 0 0 0 gpio_drive1[1]
port 100 nsew
flabel metal3 705729 134277 706005 134353 0 FreeSans 480 0 0 0 gpio_ie[1]
port 191 nsew
flabel metal3 705729 134066 706005 134142 0 FreeSans 480 0 0 0 gpio_pulldown[1]
port 305 nsew
flabel metal3 705729 133422 706005 133498 0 FreeSans 480 0 0 0 gpio_drive0[1]
port 89 nsew
flabel metal3 705729 133193 706005 133269 0 FreeSans 480 0 0 0 gpio_pullup[1]
port 343 nsew
flabel metal3 705729 132672 706005 132748 0 FreeSans 480 0 0 0 gpio_schmitt[1]
port 381 nsew
flabel metal3 705729 907706 706005 907782 0 FreeSans 480 0 0 0 gpio_ana[14]
port 466 nsew
flabel metal3 705729 821706 706005 821782 0 FreeSans 480 0 0 0 gpio_ana[13]
port 465 nsew
flabel metal3 705729 735706 706005 735782 0 FreeSans 480 0 0 0 gpio_ana[12]
port 464 nsew
flabel metal3 705729 692706 706005 692782 0 FreeSans 480 0 0 0 gpio_ana[11]
port 463 nsew
flabel metal3 705729 649706 706005 649782 0 FreeSans 480 0 0 0 gpio_ana[10]
port 462 nsew
flabel metal3 705729 606706 706005 606782 0 FreeSans 480 0 0 0 gpio_ana[9]
port 461 nsew
flabel metal3 705729 563706 706005 563782 0 FreeSans 480 0 0 0 gpio_ana[8]
port 460 nsew
flabel metal3 705729 520706 706005 520782 0 FreeSans 480 0 0 0 gpio_ana[7]
port 459 nsew
flabel metal3 705729 348706 706005 348782 0 FreeSans 480 0 0 0 gpio_ana[6]
port 458 nsew
flabel metal3 705729 305706 706005 305782 0 FreeSans 480 0 0 0 gpio_ana[5]
port 457 nsew
flabel metal3 705729 262706 706005 262782 0 FreeSans 480 0 0 0 gpio_ana[4]
port 456 nsew
flabel metal3 705729 219706 706005 219782 0 FreeSans 480 0 0 0 gpio_ana[3]
port 455 nsew
flabel metal3 705729 176706 706005 176782 0 FreeSans 480 0 0 0 gpio_ana[2]
port 454 nsew
flabel metal3 705729 90706 706005 90782 0 FreeSans 480 0 0 0 gpio_ana[0]
port 452 nsew
flabel metal3 705729 735564 706005 735640 0 FreeSans 480 0 0 0 gpio_drive1[12]
port 84 nsew
flabel metal3 705729 735422 706005 735498 0 FreeSans 480 0 0 0 gpio_drive0[12]
port 83 nsew
flabel metal3 705729 692564 706005 692640 0 FreeSans 480 0 0 0 gpio_drive1[11]
port 82 nsew
flabel metal3 705729 692422 706005 692498 0 FreeSans 480 0 0 0 gpio_drive0[11]
port 81 nsew
flabel metal3 705729 649564 706005 649640 0 FreeSans 480 0 0 0 gpio_drive1[10]
port 80 nsew
flabel metal3 705729 649422 706005 649498 0 FreeSans 480 0 0 0 gpio_drive0[10]
port 79 nsew
flabel metal3 705729 606564 706005 606640 0 FreeSans 480 0 0 0 gpio_drive1[9]
port 77 nsew
flabel metal3 705729 606422 706005 606498 0 FreeSans 480 0 0 0 gpio_drive0[9]
port 76 nsew
flabel metal3 705729 563564 706005 563640 0 FreeSans 480 0 0 0 gpio_drive1[8]
port 75 nsew
flabel metal3 705729 563422 706005 563498 0 FreeSans 480 0 0 0 gpio_drive0[8]
port 74 nsew
flabel metal3 705729 520564 706005 520640 0 FreeSans 480 0 0 0 gpio_drive1[7]
port 73 nsew
flabel metal3 705729 520422 706005 520498 0 FreeSans 480 0 0 0 gpio_drive0[7]
port 72 nsew
flabel metal3 705729 348564 706005 348640 0 FreeSans 480 0 0 0 gpio_drive1[6]
port 71 nsew
flabel metal3 705729 348422 706005 348498 0 FreeSans 480 0 0 0 gpio_drive0[6]
port 70 nsew
flabel metal3 705729 305564 706005 305640 0 FreeSans 480 0 0 0 gpio_drive1[5]
port 69 nsew
flabel metal3 705729 305422 706005 305498 0 FreeSans 480 0 0 0 gpio_drive0[5]
port 68 nsew
flabel metal3 705729 262564 706005 262640 0 FreeSans 480 0 0 0 gpio_drive1[4]
port 141 nsew
flabel metal3 705729 262422 706005 262498 0 FreeSans 480 0 0 0 gpio_drive0[4]
port 140 nsew
flabel metal3 705729 219564 706005 219640 0 FreeSans 480 0 0 0 gpio_drive1[3]
port 139 nsew
flabel metal3 705729 219422 706005 219498 0 FreeSans 480 0 0 0 gpio_drive0[3]
port 132 nsew
flabel metal3 705729 176564 706005 176640 0 FreeSans 480 0 0 0 gpio_drive1[2]
port 122 nsew
flabel metal3 705729 176422 706005 176498 0 FreeSans 480 0 0 0 gpio_drive0[2]
port 111 nsew
flabel metal3 705729 820672 706005 820748 0 FreeSans 480 0 0 0 gpio_schmitt[13]
port 374 nsew
flabel metal3 705729 821193 706005 821269 0 FreeSans 480 0 0 0 gpio_pullup[13]
port 336 nsew
flabel metal3 705729 821422 706005 821498 0 FreeSans 480 0 0 0 gpio_drive0[13]
port 85 nsew
flabel metal3 705729 821564 706005 821640 0 FreeSans 480 0 0 0 gpio_drive1[13]
port 86 nsew
flabel metal3 705729 822066 706005 822142 0 FreeSans 480 0 0 0 gpio_pulldown[13]
port 298 nsew
flabel metal3 705729 822277 706005 822353 0 FreeSans 480 0 0 0 gpio_ie[13]
port 184 nsew
flabel metal3 705729 833734 706005 833810 0 FreeSans 480 0 0 0 gpio_slew[13]
port 412 nsew
flabel metal3 705729 833880 706005 833956 0 FreeSans 480 0 0 0 gpio_out[13]
port 222 nsew
flabel metal3 705729 834026 706005 834102 0 FreeSans 480 0 0 0 gpio_oe[13]
port 260 nsew
flabel metal3 705729 834172 706005 834248 0 FreeSans 480 0 0 0 gpio_in[13]
port 146 nsew
flabel metal3 705729 734672 706005 734748 0 FreeSans 480 0 0 0 gpio_schmitt[12]
port 373 nsew
flabel metal3 705729 735193 706005 735269 0 FreeSans 480 0 0 0 gpio_pullup[12]
port 335 nsew
flabel metal3 705729 736066 706005 736142 0 FreeSans 480 0 0 0 gpio_pulldown[12]
port 297 nsew
flabel metal3 705729 736277 706005 736353 0 FreeSans 480 0 0 0 gpio_ie[12]
port 183 nsew
flabel metal3 705729 747734 706005 747810 0 FreeSans 480 0 0 0 gpio_slew[12]
port 411 nsew
flabel metal3 705729 747880 706005 747956 0 FreeSans 480 0 0 0 gpio_out[12]
port 221 nsew
flabel metal3 705729 748026 706005 748102 0 FreeSans 480 0 0 0 gpio_oe[12]
port 259 nsew
flabel metal3 705729 748172 706005 748248 0 FreeSans 480 0 0 0 gpio_in[12]
port 145 nsew
flabel metal3 705729 920172 706005 920248 0 FreeSans 480 0 0 0 gpio_in[14]
port 147 nsew
flabel metal3 705729 920026 706005 920102 0 FreeSans 480 0 0 0 gpio_oe[14]
port 261 nsew
flabel metal3 705729 919880 706005 919956 0 FreeSans 480 0 0 0 gpio_out[14]
port 223 nsew
flabel metal3 705729 919734 706005 919810 0 FreeSans 480 0 0 0 gpio_slew[14]
port 413 nsew
flabel metal3 705729 908277 706005 908353 0 FreeSans 480 0 0 0 gpio_ie[14]
port 185 nsew
flabel metal3 705729 908066 706005 908142 0 FreeSans 480 0 0 0 gpio_pulldown[14]
port 299 nsew
flabel metal3 705729 907564 706005 907640 0 FreeSans 480 0 0 0 gpio_drive1[14]
port 88 nsew
flabel metal3 705729 907422 706005 907498 0 FreeSans 480 0 0 0 gpio_drive0[14]
port 87 nsew
flabel metal3 705729 907193 706005 907269 0 FreeSans 480 0 0 0 gpio_pullup[14]
port 337 nsew
flabel metal3 705729 906672 706005 906748 0 FreeSans 480 0 0 0 gpio_schmitt[14]
port 375 nsew
flabel metal3 705729 691672 706005 691748 0 FreeSans 480 0 0 0 gpio_schmitt[11]
port 372 nsew
flabel metal3 705729 692193 706005 692269 0 FreeSans 480 0 0 0 gpio_pullup[11]
port 334 nsew
flabel metal3 705729 693066 706005 693142 0 FreeSans 480 0 0 0 gpio_pulldown[11]
port 296 nsew
flabel metal3 705729 693277 706005 693353 0 FreeSans 480 0 0 0 gpio_ie[11]
port 182 nsew
flabel metal3 705729 704734 706005 704810 0 FreeSans 480 0 0 0 gpio_slew[11]
port 410 nsew
flabel metal3 705729 704880 706005 704956 0 FreeSans 480 0 0 0 gpio_out[11]
port 220 nsew
flabel metal3 705729 705026 706005 705102 0 FreeSans 480 0 0 0 gpio_oe[11]
port 258 nsew
flabel metal3 705729 705172 706005 705248 0 FreeSans 480 0 0 0 gpio_in[11]
port 144 nsew
flabel metal3 705729 648672 706005 648748 0 FreeSans 480 0 0 0 gpio_schmitt[10]
port 371 nsew
flabel metal3 705729 649193 706005 649269 0 FreeSans 480 0 0 0 gpio_pullup[10]
port 333 nsew
flabel metal3 705729 650066 706005 650142 0 FreeSans 480 0 0 0 gpio_pulldown[10]
port 295 nsew
flabel metal3 705729 650277 706005 650353 0 FreeSans 480 0 0 0 gpio_ie[10]
port 181 nsew
flabel metal3 705729 661734 706005 661810 0 FreeSans 480 0 0 0 gpio_slew[10]
port 409 nsew
flabel metal3 705729 661880 706005 661956 0 FreeSans 480 0 0 0 gpio_out[10]
port 219 nsew
flabel metal3 705729 662026 706005 662102 0 FreeSans 480 0 0 0 gpio_oe[10]
port 257 nsew
flabel metal3 705729 662172 706005 662248 0 FreeSans 480 0 0 0 gpio_in[10]
port 143 nsew
flabel metal3 705729 605672 706005 605748 0 FreeSans 480 0 0 0 gpio_schmitt[9]
port 407 nsew
flabel metal3 705729 606193 706005 606269 0 FreeSans 480 0 0 0 gpio_pullup[9]
port 369 nsew
flabel metal3 705729 607066 706005 607142 0 FreeSans 480 0 0 0 gpio_pulldown[9]
port 331 nsew
flabel metal3 705729 607277 706005 607353 0 FreeSans 480 0 0 0 gpio_ie[9]
port 217 nsew
flabel metal3 705729 618734 706005 618810 0 FreeSans 480 0 0 0 gpio_slew[9]
port 445 nsew
flabel metal3 705729 618880 706005 618956 0 FreeSans 480 0 0 0 gpio_out[9]
port 255 nsew
flabel metal3 705729 619026 706005 619102 0 FreeSans 480 0 0 0 gpio_oe[9]
port 293 nsew
flabel metal3 705729 619172 706005 619248 0 FreeSans 480 0 0 0 gpio_in[9]
port 179 nsew
flabel metal3 705729 562672 706005 562748 0 FreeSans 480 0 0 0 gpio_schmitt[8]
port 406 nsew
flabel metal3 705729 563193 706005 563269 0 FreeSans 480 0 0 0 gpio_pullup[8]
port 368 nsew
flabel metal3 705729 564066 706005 564142 0 FreeSans 480 0 0 0 gpio_pulldown[8]
port 330 nsew
flabel metal3 705729 564277 706005 564353 0 FreeSans 480 0 0 0 gpio_ie[8]
port 216 nsew
flabel metal3 705729 575734 706005 575810 0 FreeSans 480 0 0 0 gpio_slew[8]
port 444 nsew
flabel metal3 705729 575880 706005 575956 0 FreeSans 480 0 0 0 gpio_out[8]
port 254 nsew
flabel metal3 705729 576026 706005 576102 0 FreeSans 480 0 0 0 gpio_oe[8]
port 292 nsew
flabel metal3 705729 576172 706005 576248 0 FreeSans 480 0 0 0 gpio_in[8]
port 178 nsew
flabel metal3 705729 519672 706005 519748 0 FreeSans 480 0 0 0 gpio_schmitt[7]
port 405 nsew
flabel metal3 705729 520193 706005 520269 0 FreeSans 480 0 0 0 gpio_pullup[7]
port 367 nsew
flabel metal3 705729 521066 706005 521142 0 FreeSans 480 0 0 0 gpio_pulldown[7]
port 329 nsew
flabel metal3 705729 521277 706005 521353 0 FreeSans 480 0 0 0 gpio_ie[7]
port 215 nsew
flabel metal3 705729 532734 706005 532810 0 FreeSans 480 0 0 0 gpio_slew[7]
port 443 nsew
flabel metal3 705729 532880 706005 532956 0 FreeSans 480 0 0 0 gpio_out[7]
port 253 nsew
flabel metal3 705729 533026 706005 533102 0 FreeSans 480 0 0 0 gpio_oe[7]
port 291 nsew
flabel metal3 705729 533172 706005 533248 0 FreeSans 480 0 0 0 gpio_in[7]
port 177 nsew
flabel metal3 705729 347672 706005 347748 0 FreeSans 480 0 0 0 gpio_schmitt[6]
port 404 nsew
flabel metal3 705729 348193 706005 348269 0 FreeSans 480 0 0 0 gpio_pullup[6]
port 366 nsew
flabel metal3 705729 349066 706005 349142 0 FreeSans 480 0 0 0 gpio_pulldown[6]
port 328 nsew
flabel metal3 705729 349277 706005 349353 0 FreeSans 480 0 0 0 gpio_ie[6]
port 214 nsew
flabel metal3 705729 360734 706005 360810 0 FreeSans 480 0 0 0 gpio_slew[6]
port 442 nsew
flabel metal3 705729 360880 706005 360956 0 FreeSans 480 0 0 0 gpio_out[6]
port 252 nsew
flabel metal3 705729 361026 706005 361102 0 FreeSans 480 0 0 0 gpio_oe[6]
port 290 nsew
flabel metal3 705729 361172 706005 361248 0 FreeSans 480 0 0 0 gpio_in[6]
port 176 nsew
flabel metal3 705729 304672 706005 304748 0 FreeSans 480 0 0 0 gpio_schmitt[5]
port 403 nsew
flabel metal3 705729 305193 706005 305269 0 FreeSans 480 0 0 0 gpio_pullup[5]
port 365 nsew
flabel metal3 705729 306066 706005 306142 0 FreeSans 480 0 0 0 gpio_pulldown[5]
port 327 nsew
flabel metal3 705729 306277 706005 306353 0 FreeSans 480 0 0 0 gpio_ie[5]
port 213 nsew
flabel metal3 705729 317734 706005 317810 0 FreeSans 480 0 0 0 gpio_slew[5]
port 441 nsew
flabel metal3 705729 317880 706005 317956 0 FreeSans 480 0 0 0 gpio_out[5]
port 251 nsew
flabel metal3 705729 318026 706005 318102 0 FreeSans 480 0 0 0 gpio_oe[5]
port 289 nsew
flabel metal3 705729 318172 706005 318248 0 FreeSans 480 0 0 0 gpio_in[5]
port 175 nsew
flabel metal3 705729 261672 706005 261748 0 FreeSans 480 0 0 0 gpio_schmitt[4]
port 402 nsew
flabel metal3 705729 262193 706005 262269 0 FreeSans 480 0 0 0 gpio_pullup[4]
port 364 nsew
flabel metal3 705729 263066 706005 263142 0 FreeSans 480 0 0 0 gpio_pulldown[4]
port 326 nsew
flabel metal3 705729 263277 706005 263353 0 FreeSans 480 0 0 0 gpio_ie[4]
port 212 nsew
flabel metal3 705729 274734 706005 274810 0 FreeSans 480 0 0 0 gpio_slew[4]
port 440 nsew
flabel metal3 705729 274880 706005 274956 0 FreeSans 480 0 0 0 gpio_out[4]
port 250 nsew
flabel metal3 705729 275026 706005 275102 0 FreeSans 480 0 0 0 gpio_oe[4]
port 288 nsew
flabel metal3 705729 275172 706005 275248 0 FreeSans 480 0 0 0 gpio_in[4]
port 174 nsew
flabel metal3 705729 218672 706005 218748 0 FreeSans 480 0 0 0 gpio_schmitt[3]
port 401 nsew
flabel metal3 705729 219193 706005 219269 0 FreeSans 480 0 0 0 gpio_pullup[3]
port 363 nsew
flabel metal3 705729 220066 706005 220142 0 FreeSans 480 0 0 0 gpio_pulldown[3]
port 325 nsew
flabel metal3 705729 220277 706005 220353 0 FreeSans 480 0 0 0 gpio_ie[3]
port 211 nsew
flabel metal3 705729 231734 706005 231810 0 FreeSans 480 0 0 0 gpio_slew[3]
port 439 nsew
flabel metal3 705729 231880 706005 231956 0 FreeSans 480 0 0 0 gpio_out[3]
port 249 nsew
flabel metal3 705729 232026 706005 232102 0 FreeSans 480 0 0 0 gpio_oe[3]
port 287 nsew
flabel metal3 705729 232172 706005 232248 0 FreeSans 480 0 0 0 gpio_in[3]
port 173 nsew
flabel metal3 705729 175672 706005 175748 0 FreeSans 480 0 0 0 gpio_schmitt[2]
port 392 nsew
flabel metal3 705729 176193 706005 176269 0 FreeSans 480 0 0 0 gpio_pullup[2]
port 354 nsew
flabel metal3 705729 177066 706005 177142 0 FreeSans 480 0 0 0 gpio_pulldown[2]
port 316 nsew
flabel metal3 705729 177277 706005 177353 0 FreeSans 480 0 0 0 gpio_ie[2]
port 202 nsew
flabel metal3 705729 188734 706005 188810 0 FreeSans 480 0 0 0 gpio_slew[2]
port 430 nsew
flabel metal3 705729 188880 706005 188956 0 FreeSans 480 0 0 0 gpio_out[2]
port 240 nsew
flabel metal3 705729 189026 706005 189102 0 FreeSans 480 0 0 0 gpio_oe[2]
port 278 nsew
flabel metal3 705729 189172 706005 189248 0 FreeSans 480 0 0 0 gpio_in[2]
port 164 nsew
flabel metal3 705729 103172 706005 103248 0 FreeSans 480 0 0 0 gpio_in[0]
port 142 nsew
flabel metal3 705729 103026 706005 103102 0 FreeSans 480 0 0 0 gpio_oe[0]
port 256 nsew
flabel metal3 705729 102880 706005 102956 0 FreeSans 480 0 0 0 gpio_out[0]
port 218 nsew
flabel metal3 705729 102734 706005 102810 0 FreeSans 480 0 0 0 gpio_slew[0]
port 408 nsew
flabel metal3 705729 91277 706005 91353 0 FreeSans 480 0 0 0 gpio_ie[0]
port 180 nsew
flabel metal3 705729 91066 706005 91142 0 FreeSans 480 0 0 0 gpio_pulldown[0]
port 294 nsew
flabel metal3 705729 90564 706005 90640 0 FreeSans 480 0 0 0 gpio_drive1[0]
port 78 nsew
flabel metal3 705729 90422 706005 90498 0 FreeSans 480 0 0 0 gpio_drive0[0]
port 67 nsew
flabel metal3 705729 90193 706005 90269 0 FreeSans 480 0 0 0 gpio_pullup[0]
port 332 nsew
flabel metal3 705729 89672 706005 89748 0 FreeSans 480 0 0 0 gpio_schmitt[0]
port 370 nsew
flabel metal3 69995 167752 70271 167828 0 FreeSans 480 180 0 0 gpio_in[37]
port 172 nsew
flabel metal3 69995 167898 70271 167974 0 FreeSans 480 180 0 0 gpio_oe[37]
port 286 nsew
flabel metal3 69995 168044 70271 168120 0 FreeSans 480 180 0 0 gpio_out[37]
port 248 nsew
flabel metal3 69995 168190 70271 168266 0 FreeSans 480 180 0 0 gpio_slew[37]
port 438 nsew
flabel metal3 69995 179647 70271 179723 0 FreeSans 480 180 0 0 gpio_ie[37]
port 210 nsew
flabel metal3 69995 179858 70271 179934 0 FreeSans 480 180 0 0 gpio_pulldown[37]
port 324 nsew
flabel metal3 69995 180360 70271 180436 0 FreeSans 480 180 0 0 gpio_drive1[37]
port 138 nsew
flabel metal3 69995 180502 70271 180578 0 FreeSans 480 180 0 0 gpio_drive0[37]
port 137 nsew
flabel metal3 69995 180731 70271 180807 0 FreeSans 480 180 0 0 gpio_pullup[37]
port 362 nsew
flabel metal3 69995 181252 70271 181328 0 FreeSans 480 180 0 0 gpio_schmitt[37]
port 400 nsew
flabel metal3 69995 208752 70271 208828 0 FreeSans 480 180 0 0 gpio_in[36]
port 171 nsew
flabel metal3 69995 208898 70271 208974 0 FreeSans 480 180 0 0 gpio_oe[36]
port 285 nsew
flabel metal3 69995 209044 70271 209120 0 FreeSans 480 180 0 0 gpio_out[36]
port 247 nsew
flabel metal3 69995 209190 70271 209266 0 FreeSans 480 180 0 0 gpio_slew[36]
port 437 nsew
flabel metal3 69995 220647 70271 220723 0 FreeSans 480 180 0 0 gpio_ie[36]
port 209 nsew
flabel metal3 69995 220858 70271 220934 0 FreeSans 480 180 0 0 gpio_pulldown[36]
port 323 nsew
flabel metal3 69995 221360 70271 221436 0 FreeSans 480 180 0 0 gpio_drive1[36]
port 136 nsew
flabel metal3 69995 221502 70271 221578 0 FreeSans 480 180 0 0 gpio_drive0[36]
port 135 nsew
flabel metal3 69995 221731 70271 221807 0 FreeSans 480 180 0 0 gpio_pullup[36]
port 361 nsew
flabel metal3 69995 222252 70271 222328 0 FreeSans 480 180 0 0 gpio_schmitt[36]
port 399 nsew
flabel metal3 69995 249752 70271 249828 0 FreeSans 480 180 0 0 gpio_in[35]
port 170 nsew
flabel metal3 69995 249898 70271 249974 0 FreeSans 480 180 0 0 gpio_oe[35]
port 284 nsew
flabel metal3 69995 250044 70271 250120 0 FreeSans 480 180 0 0 gpio_out[35]
port 246 nsew
flabel metal3 69995 250190 70271 250266 0 FreeSans 480 180 0 0 gpio_slew[35]
port 436 nsew
flabel metal3 69995 261647 70271 261723 0 FreeSans 480 180 0 0 gpio_ie[35]
port 208 nsew
flabel metal3 69995 261858 70271 261934 0 FreeSans 480 180 0 0 gpio_pulldown[35]
port 322 nsew
flabel metal3 69995 262360 70271 262436 0 FreeSans 480 180 0 0 gpio_drive1[35]
port 134 nsew
flabel metal3 69995 262502 70271 262578 0 FreeSans 480 180 0 0 gpio_drive0[35]
port 133 nsew
flabel metal3 69995 262731 70271 262807 0 FreeSans 480 180 0 0 gpio_pullup[35]
port 360 nsew
flabel metal3 69995 263252 70271 263328 0 FreeSans 480 180 0 0 gpio_schmitt[35]
port 398 nsew
flabel metal3 69995 290752 70271 290828 0 FreeSans 480 180 0 0 gpio_in[34]
port 169 nsew
flabel metal3 69995 262218 70271 262294 0 FreeSans 480 180 0 0 gpio_ana[35]
port 487 nsew
flabel metal3 69995 221218 70271 221294 0 FreeSans 480 180 0 0 gpio_ana[36]
port 488 nsew
flabel metal3 69995 180218 70271 180294 0 FreeSans 480 180 0 0 gpio_ana[37]
port 489 nsew
flabel metal3 69971 289178 70271 289254 0 FreeSans 480 0 0 0 gpio_loopback_zero[34]
port 564 nsew
flabel metal3 69971 207178 70271 207254 0 FreeSans 480 0 0 0 gpio_loopback_zero[36]
port 568 nsew
flabel metal3 69971 371178 70271 371254 0 FreeSans 480 0 0 0 gpio_loopback_zero[32]
port 560 nsew
flabel metal3 69971 535366 70271 535442 0 FreeSans 480 0 0 0 gpio_loopback_one[30]
port 557 nsew
flabel metal3 69971 535178 70271 535254 0 FreeSans 480 0 0 0 gpio_loopback_zero[30]
port 556 nsew
flabel metal3 69971 617366 70271 617442 0 FreeSans 480 0 0 0 gpio_loopback_one[28]
port 553 nsew
flabel metal3 69971 617178 70271 617254 0 FreeSans 480 0 0 0 gpio_loopback_zero[28]
port 552 nsew
flabel metal3 69971 699366 70271 699442 0 FreeSans 480 0 0 0 gpio_loopback_one[26]
port 549 nsew
flabel metal3 69971 699178 70271 699254 0 FreeSans 480 0 0 0 gpio_loopback_zero[26]
port 548 nsew
flabel metal3 69971 904366 70271 904442 0 FreeSans 480 0 0 0 gpio_loopback_one[24]
port 545 nsew
flabel metal3 69995 303218 70271 303294 0 FreeSans 480 180 0 0 gpio_ana[34]
port 486 nsew
flabel metal3 69995 344218 70271 344294 0 FreeSans 480 180 0 0 gpio_ana[33]
port 485 nsew
flabel metal3 69995 385218 70271 385294 0 FreeSans 480 180 0 0 gpio_ana[32]
port 484 nsew
flabel metal3 69995 508218 70271 508294 0 FreeSans 480 180 0 0 gpio_ana[31]
port 483 nsew
flabel metal3 69995 549218 70271 549294 0 FreeSans 480 180 0 0 gpio_ana[30]
port 482 nsew
flabel metal3 69995 590218 70271 590294 0 FreeSans 480 180 0 0 gpio_ana[29]
port 481 nsew
flabel metal3 69995 631218 70271 631294 0 FreeSans 480 180 0 0 gpio_ana[28]
port 480 nsew
flabel metal3 69995 672218 70271 672294 0 FreeSans 480 180 0 0 gpio_ana[27]
port 479 nsew
flabel metal3 69995 713218 70271 713294 0 FreeSans 480 180 0 0 gpio_ana[26]
port 478 nsew
flabel metal3 69995 754218 70271 754294 0 FreeSans 480 180 0 0 gpio_ana[25]
port 477 nsew
flabel metal3 69995 918218 70271 918294 0 FreeSans 480 180 0 0 gpio_ana[24]
port 476 nsew
flabel metal3 69995 549502 70271 549578 0 FreeSans 480 180 0 0 gpio_drive0[30]
port 66 nsew
flabel metal3 69995 549360 70271 549436 0 FreeSans 480 180 0 0 gpio_drive1[30]
port 123 nsew
flabel metal3 69995 919252 70271 919328 0 FreeSans 480 180 0 0 gpio_schmitt[24]
port 386 nsew
flabel metal3 69995 918731 70271 918807 0 FreeSans 480 180 0 0 gpio_pullup[24]
port 348 nsew
flabel metal3 69995 918502 70271 918578 0 FreeSans 480 180 0 0 gpio_drive0[24]
port 109 nsew
flabel metal3 69995 918360 70271 918436 0 FreeSans 480 180 0 0 gpio_drive1[24]
port 110 nsew
flabel metal3 69995 917858 70271 917934 0 FreeSans 480 180 0 0 gpio_pulldown[24]
port 310 nsew
flabel metal3 69995 917647 70271 917723 0 FreeSans 480 180 0 0 gpio_ie[24]
port 196 nsew
flabel metal3 69995 906190 70271 906266 0 FreeSans 480 180 0 0 gpio_slew[24]
port 424 nsew
flabel metal3 69995 906044 70271 906120 0 FreeSans 480 180 0 0 gpio_out[24]
port 234 nsew
flabel metal3 69995 905898 70271 905974 0 FreeSans 480 180 0 0 gpio_oe[24]
port 272 nsew
flabel metal3 69995 905752 70271 905828 0 FreeSans 480 180 0 0 gpio_in[24]
port 158 nsew
flabel metal3 69995 755252 70271 755328 0 FreeSans 480 180 0 0 gpio_schmitt[25]
port 387 nsew
flabel metal3 69995 754731 70271 754807 0 FreeSans 480 180 0 0 gpio_pullup[25]
port 349 nsew
flabel metal3 69995 754502 70271 754578 0 FreeSans 480 180 0 0 gpio_drive0[25]
port 113 nsew
flabel metal3 69995 754360 70271 754436 0 FreeSans 480 180 0 0 gpio_drive1[25]
port 112 nsew
flabel metal3 69995 753858 70271 753934 0 FreeSans 480 180 0 0 gpio_pulldown[25]
port 311 nsew
flabel metal3 69995 753647 70271 753723 0 FreeSans 480 180 0 0 gpio_ie[25]
port 197 nsew
flabel metal3 69995 742190 70271 742266 0 FreeSans 480 180 0 0 gpio_slew[25]
port 425 nsew
flabel metal3 69995 742044 70271 742120 0 FreeSans 480 180 0 0 gpio_out[25]
port 235 nsew
flabel metal3 69995 741898 70271 741974 0 FreeSans 480 180 0 0 gpio_oe[25]
port 273 nsew
flabel metal3 69995 741752 70271 741828 0 FreeSans 480 180 0 0 gpio_in[25]
port 159 nsew
flabel metal3 69995 714252 70271 714328 0 FreeSans 480 180 0 0 gpio_schmitt[26]
port 388 nsew
flabel metal3 69995 713731 70271 713807 0 FreeSans 480 180 0 0 gpio_pullup[26]
port 350 nsew
flabel metal3 69995 713502 70271 713578 0 FreeSans 480 180 0 0 gpio_drive0[26]
port 114 nsew
flabel metal3 69995 713360 70271 713436 0 FreeSans 480 180 0 0 gpio_drive1[26]
port 115 nsew
flabel metal3 69995 712858 70271 712934 0 FreeSans 480 180 0 0 gpio_pulldown[26]
port 312 nsew
flabel metal3 69995 712647 70271 712723 0 FreeSans 480 180 0 0 gpio_ie[26]
port 198 nsew
flabel metal3 69995 701190 70271 701266 0 FreeSans 480 180 0 0 gpio_slew[26]
port 426 nsew
flabel metal3 69995 701044 70271 701120 0 FreeSans 480 180 0 0 gpio_out[26]
port 236 nsew
flabel metal3 69995 700898 70271 700974 0 FreeSans 480 180 0 0 gpio_oe[26]
port 274 nsew
flabel metal3 69995 700752 70271 700828 0 FreeSans 480 180 0 0 gpio_in[26]
port 160 nsew
flabel metal3 69995 673252 70271 673328 0 FreeSans 480 180 0 0 gpio_schmitt[27]
port 389 nsew
flabel metal3 69995 672731 70271 672807 0 FreeSans 480 180 0 0 gpio_pullup[27]
port 351 nsew
flabel metal3 69995 672502 70271 672578 0 FreeSans 480 180 0 0 gpio_drive0[27]
port 116 nsew
flabel metal3 69995 672360 70271 672436 0 FreeSans 480 180 0 0 gpio_drive1[27]
port 117 nsew
flabel metal3 69995 671858 70271 671934 0 FreeSans 480 180 0 0 gpio_pulldown[27]
port 313 nsew
flabel metal3 69995 671647 70271 671723 0 FreeSans 480 180 0 0 gpio_ie[27]
port 199 nsew
flabel metal3 69995 660190 70271 660266 0 FreeSans 480 180 0 0 gpio_slew[27]
port 427 nsew
flabel metal3 69995 660044 70271 660120 0 FreeSans 480 180 0 0 gpio_out[27]
port 237 nsew
flabel metal3 69995 659898 70271 659974 0 FreeSans 480 180 0 0 gpio_oe[27]
port 275 nsew
flabel metal3 69995 659752 70271 659828 0 FreeSans 480 180 0 0 gpio_in[27]
port 161 nsew
flabel metal3 69995 632252 70271 632328 0 FreeSans 480 180 0 0 gpio_schmitt[28]
port 390 nsew
flabel metal3 69995 631731 70271 631807 0 FreeSans 480 180 0 0 gpio_pullup[28]
port 352 nsew
flabel metal3 69995 631502 70271 631578 0 FreeSans 480 180 0 0 gpio_drive0[28]
port 118 nsew
flabel metal3 69995 631360 70271 631436 0 FreeSans 480 180 0 0 gpio_drive1[28]
port 119 nsew
flabel metal3 69995 630858 70271 630934 0 FreeSans 480 180 0 0 gpio_pulldown[28]
port 314 nsew
flabel metal3 69995 630647 70271 630723 0 FreeSans 480 180 0 0 gpio_ie[28]
port 200 nsew
flabel metal3 69995 619190 70271 619266 0 FreeSans 480 180 0 0 gpio_slew[28]
port 428 nsew
flabel metal3 69995 619044 70271 619120 0 FreeSans 480 180 0 0 gpio_out[28]
port 238 nsew
flabel metal3 69995 618898 70271 618974 0 FreeSans 480 180 0 0 gpio_oe[28]
port 276 nsew
flabel metal3 69995 618752 70271 618828 0 FreeSans 480 180 0 0 gpio_in[28]
port 162 nsew
flabel metal3 69995 591252 70271 591328 0 FreeSans 480 180 0 0 gpio_schmitt[29]
port 391 nsew
flabel metal3 69995 590731 70271 590807 0 FreeSans 480 180 0 0 gpio_pullup[29]
port 353 nsew
flabel metal3 69995 590502 70271 590578 0 FreeSans 480 180 0 0 gpio_drive0[29]
port 120 nsew
flabel metal3 69995 590360 70271 590436 0 FreeSans 480 180 0 0 gpio_drive1[29]
port 121 nsew
flabel metal3 69995 589858 70271 589934 0 FreeSans 480 180 0 0 gpio_pulldown[29]
port 315 nsew
flabel metal3 69995 589647 70271 589723 0 FreeSans 480 180 0 0 gpio_ie[29]
port 201 nsew
flabel metal3 69995 578190 70271 578266 0 FreeSans 480 180 0 0 gpio_slew[29]
port 429 nsew
flabel metal3 69995 578044 70271 578120 0 FreeSans 480 180 0 0 gpio_out[29]
port 239 nsew
flabel metal3 69995 577898 70271 577974 0 FreeSans 480 180 0 0 gpio_oe[29]
port 277 nsew
flabel metal3 69995 577752 70271 577828 0 FreeSans 480 180 0 0 gpio_in[29]
port 163 nsew
flabel metal3 69995 550252 70271 550328 0 FreeSans 480 180 0 0 gpio_schmitt[30]
port 393 nsew
flabel metal3 69995 549731 70271 549807 0 FreeSans 480 180 0 0 gpio_pullup[30]
port 355 nsew
flabel metal3 69995 548858 70271 548934 0 FreeSans 480 180 0 0 gpio_pulldown[30]
port 317 nsew
flabel metal3 69995 548647 70271 548723 0 FreeSans 480 180 0 0 gpio_ie[30]
port 203 nsew
flabel metal3 69995 537190 70271 537266 0 FreeSans 480 180 0 0 gpio_slew[30]
port 431 nsew
flabel metal3 69995 537044 70271 537120 0 FreeSans 480 180 0 0 gpio_out[30]
port 241 nsew
flabel metal3 69995 536898 70271 536974 0 FreeSans 480 180 0 0 gpio_oe[30]
port 279 nsew
flabel metal3 69995 536752 70271 536828 0 FreeSans 480 180 0 0 gpio_in[30]
port 165 nsew
flabel metal3 69995 509252 70271 509328 0 FreeSans 480 180 0 0 gpio_schmitt[31]
port 394 nsew
flabel metal3 69995 508731 70271 508807 0 FreeSans 480 180 0 0 gpio_pullup[31]
port 356 nsew
flabel metal3 69995 508502 70271 508578 0 FreeSans 480 180 0 0 gpio_drive0[31]
port 124 nsew
flabel metal3 69995 508360 70271 508436 0 FreeSans 480 180 0 0 gpio_drive1[31]
port 125 nsew
flabel metal3 69995 507858 70271 507934 0 FreeSans 480 180 0 0 gpio_pulldown[31]
port 318 nsew
flabel metal3 69995 507647 70271 507723 0 FreeSans 480 180 0 0 gpio_ie[31]
port 204 nsew
flabel metal3 69995 496190 70271 496266 0 FreeSans 480 180 0 0 gpio_slew[31]
port 432 nsew
flabel metal3 69995 496044 70271 496120 0 FreeSans 480 180 0 0 gpio_out[31]
port 242 nsew
flabel metal3 69995 495898 70271 495974 0 FreeSans 480 180 0 0 gpio_oe[31]
port 280 nsew
flabel metal3 69995 495752 70271 495828 0 FreeSans 480 180 0 0 gpio_in[31]
port 166 nsew
flabel metal3 69995 386252 70271 386328 0 FreeSans 480 180 0 0 gpio_schmitt[32]
port 395 nsew
flabel metal3 69995 385731 70271 385807 0 FreeSans 480 180 0 0 gpio_pullup[32]
port 357 nsew
flabel metal3 69995 385502 70271 385578 0 FreeSans 480 180 0 0 gpio_drive0[32]
port 126 nsew
flabel metal3 69995 385360 70271 385436 0 FreeSans 480 180 0 0 gpio_drive1[32]
port 127 nsew
flabel metal3 69995 384858 70271 384934 0 FreeSans 480 180 0 0 gpio_pulldown[32]
port 319 nsew
flabel metal3 69995 384647 70271 384723 0 FreeSans 480 180 0 0 gpio_ie[32]
port 205 nsew
flabel metal3 69995 373190 70271 373266 0 FreeSans 480 180 0 0 gpio_slew[32]
port 433 nsew
flabel metal3 69995 373044 70271 373120 0 FreeSans 480 180 0 0 gpio_out[32]
port 243 nsew
flabel metal3 69995 372898 70271 372974 0 FreeSans 480 180 0 0 gpio_oe[32]
port 281 nsew
flabel metal3 69995 372752 70271 372828 0 FreeSans 480 180 0 0 gpio_in[32]
port 167 nsew
flabel metal3 69995 345252 70271 345328 0 FreeSans 480 180 0 0 gpio_schmitt[33]
port 396 nsew
flabel metal3 69995 344731 70271 344807 0 FreeSans 480 180 0 0 gpio_pullup[33]
port 358 nsew
flabel metal3 69995 344502 70271 344578 0 FreeSans 480 180 0 0 gpio_drive0[33]
port 128 nsew
flabel metal3 69995 344360 70271 344436 0 FreeSans 480 180 0 0 gpio_drive1[33]
port 129 nsew
flabel metal3 69995 343858 70271 343934 0 FreeSans 480 180 0 0 gpio_pulldown[33]
port 320 nsew
flabel metal3 69995 343647 70271 343723 0 FreeSans 480 180 0 0 gpio_ie[33]
port 206 nsew
flabel metal3 69995 332190 70271 332266 0 FreeSans 480 180 0 0 gpio_slew[33]
port 434 nsew
flabel metal3 69995 332044 70271 332120 0 FreeSans 480 180 0 0 gpio_out[33]
port 244 nsew
flabel metal3 69995 331898 70271 331974 0 FreeSans 480 180 0 0 gpio_oe[33]
port 282 nsew
flabel metal3 69995 331752 70271 331828 0 FreeSans 480 180 0 0 gpio_in[33]
port 168 nsew
flabel metal3 69995 304252 70271 304328 0 FreeSans 480 180 0 0 gpio_schmitt[34]
port 397 nsew
flabel metal3 69995 303731 70271 303807 0 FreeSans 480 180 0 0 gpio_pullup[34]
port 359 nsew
flabel metal3 69995 303502 70271 303578 0 FreeSans 480 180 0 0 gpio_drive0[34]
port 130 nsew
flabel metal3 69995 303360 70271 303436 0 FreeSans 480 180 0 0 gpio_drive1[34]
port 131 nsew
flabel metal3 69995 302858 70271 302934 0 FreeSans 480 180 0 0 gpio_pulldown[34]
port 321 nsew
flabel metal3 69995 302647 70271 302723 0 FreeSans 480 180 0 0 gpio_ie[34]
port 207 nsew
flabel metal3 69995 291190 70271 291266 0 FreeSans 480 180 0 0 gpio_slew[34]
port 435 nsew
flabel metal3 69995 291044 70271 291120 0 FreeSans 480 180 0 0 gpio_out[34]
port 245 nsew
flabel metal3 69995 290898 70271 290974 0 FreeSans 480 180 0 0 gpio_oe[34]
port 283 nsew
flabel metal2 590707 69900 590783 70200 0 FreeSans 480 90 0 0 por_h
port 589 nsew
flabel metal2 591290 69900 591366 70200 0 FreeSans 480 90 0 0 porb_h
port 590 nsew
flabel metal2 593218 69900 593294 70200 0 FreeSans 480 90 0 0 porb_l
port 591 nsew
flabel metal2 507707 69900 507783 70200 0 FreeSans 480 90 0 0 mask_rev[0]
port 592 nsew
flabel metal2 508290 69900 508366 70200 0 FreeSans 480 90 0 0 mask_rev[1]
port 593 nsew
flabel metal2 509707 69900 509783 70200 0 FreeSans 480 90 0 0 mask_rev[2]
port 594 nsew
flabel metal2 510290 69900 510366 70200 0 FreeSans 480 90 0 0 mask_rev[3]
port 595 nsew
flabel metal2 511707 69900 511783 70200 0 FreeSans 480 90 0 0 mask_rev[4]
port 596 nsew
flabel metal2 512290 69900 512366 70200 0 FreeSans 480 90 0 0 mask_rev[5]
port 597 nsew
flabel metal2 513707 69900 513783 70200 0 FreeSans 480 90 0 0 mask_rev[6]
port 598 nsew
flabel metal2 514290 69900 514366 70200 0 FreeSans 480 90 0 0 mask_rev[7]
port 599 nsew
flabel metal2 515707 69900 515783 70200 0 FreeSans 480 90 0 0 mask_rev[8]
port 600 nsew
flabel metal2 516290 69900 516366 70200 0 FreeSans 480 90 0 0 mask_rev[9]
port 601 nsew
flabel metal2 517707 69900 517783 70200 0 FreeSans 480 90 0 0 mask_rev[10]
port 602 nsew
flabel metal2 518290 69900 518366 70200 0 FreeSans 480 90 0 0 mask_rev[11]
port 603 nsew
flabel metal2 519707 69900 519783 70200 0 FreeSans 480 90 0 0 mask_rev[12]
port 604 nsew
flabel metal2 520290 69900 520366 70200 0 FreeSans 480 90 0 0 mask_rev[13]
port 605 nsew
flabel metal2 521707 69900 521783 70200 0 FreeSans 480 90 0 0 mask_rev[14]
port 606 nsew
flabel metal2 522290 69900 522366 70200 0 FreeSans 480 90 0 0 mask_rev[15]
port 607 nsew
flabel metal2 523707 69900 523783 70200 0 FreeSans 480 90 0 0 mask_rev[16]
port 608 nsew
flabel metal2 524290 69900 524366 70200 0 FreeSans 480 90 0 0 mask_rev[17]
port 609 nsew
flabel metal2 525707 69900 525783 70200 0 FreeSans 480 90 0 0 mask_rev[18]
port 610 nsew
flabel metal2 526290 69900 526366 70200 0 FreeSans 480 90 0 0 mask_rev[19]
port 611 nsew
flabel metal2 527707 69900 527783 70200 0 FreeSans 480 90 0 0 mask_rev[20]
port 612 nsew
flabel metal2 528290 69900 528366 70200 0 FreeSans 480 90 0 0 mask_rev[21]
port 613 nsew
flabel metal2 529707 69900 529783 70200 0 FreeSans 480 90 0 0 mask_rev[22]
port 614 nsew
flabel metal2 530290 69900 530366 70200 0 FreeSans 480 90 0 0 mask_rev[23]
port 615 nsew
flabel metal2 531707 69900 531783 70200 0 FreeSans 480 90 0 0 mask_rev[24]
port 616 nsew
flabel metal2 532290 69900 532366 70200 0 FreeSans 480 90 0 0 mask_rev[25]
port 617 nsew
flabel metal2 533707 69900 533783 70200 0 FreeSans 480 90 0 0 mask_rev[26]
port 618 nsew
flabel metal2 534290 69900 534366 70200 0 FreeSans 480 90 0 0 mask_rev[27]
port 619 nsew
flabel metal2 535707 69900 535783 70200 0 FreeSans 480 90 0 0 mask_rev[28]
port 620 nsew
flabel metal2 536290 69900 536366 70200 0 FreeSans 480 90 0 0 mask_rev[29]
port 621 nsew
flabel metal2 537707 69900 537783 70200 0 FreeSans 480 90 0 0 mask_rev[30]
port 622 nsew
flabel metal2 538290 69900 538366 70200 0 FreeSans 480 90 0 0 mask_rev[31]
port 623 nsew
flabel metal2 159178 69900 159254 70200 0 FreeSans 480 90 0 0 resetb_loopback_zero
port 588 nsew
flabel metal2 159366 69900 159442 70200 0 FreeSans 480 90 0 0 resetb_loopback_one
port 587 nsew
flabel metal4 105272 70000 107172 70200 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 107752 70000 109802 70200 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 110122 70000 112172 70200 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 112828 70000 114878 70200 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 115198 70000 117248 70200 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 117828 70000 119728 70200 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 270272 70000 272172 70200 0 FreeSans 1600 0 0 0 vssd
port 625 nsew
flabel metal4 272752 70000 274802 70200 0 FreeSans 1600 0 0 0 vssd
port 625 nsew
flabel metal4 275122 70000 277172 70200 0 FreeSans 1600 0 0 0 vssd
port 625 nsew
flabel metal4 277828 70000 279878 70200 0 FreeSans 1600 0 0 0 vssd
port 625 nsew
flabel metal4 280198 70000 282248 70200 0 FreeSans 1600 0 0 0 vssd
port 625 nsew
flabel metal4 282828 70000 284728 70200 0 FreeSans 1600 0 0 0 vssd
port 625 nsew
flabel metal4 600272 70000 602172 70200 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 602752 70000 604802 70200 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 605122 70000 607172 70200 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 607828 70000 609878 70200 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 610198 70000 612248 70200 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 612828 70000 614728 70200 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 655272 69999 657172 70199 0 FreeSans 1600 0 0 0 vddio
port 626 nsew
flabel metal4 657752 69999 659802 70199 0 FreeSans 1600 0 0 0 vddio
port 626 nsew
flabel metal4 660122 69999 662172 70199 0 FreeSans 1600 0 0 0 vddio
port 626 nsew
flabel metal4 662828 69999 664878 70199 0 FreeSans 1600 0 0 0 vddio
port 626 nsew
flabel metal4 665198 69999 667248 70199 0 FreeSans 1600 0 0 0 vddio
port 626 nsew
flabel metal4 667828 69999 669728 70199 0 FreeSans 1600 0 0 0 vddio
port 626 nsew
flabel metal4 379272 943800 381172 944000 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 381752 943800 383802 944000 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 384122 943800 386172 944000 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 386828 943800 388878 944000 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 389198 943800 391248 944000 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 391828 943800 393728 944000 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 599272 943800 601172 944000 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 601752 943800 603802 944000 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 604122 943800 606172 944000 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 606828 943800 608878 944000 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 609198 943800 611248 944000 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal4 611828 943800 613728 944000 0 FreeSans 1600 0 0 0 vssio
port 624 nsew
flabel metal5 705730 390272 706000 392172 0 FreeSans 1600 90 0 0 vssio
port 624 nsew
flabel metal5 705730 392752 706000 394802 0 FreeSans 1600 90 0 0 vssio
port 624 nsew
flabel metal5 705730 395122 706000 397172 0 FreeSans 1600 90 0 0 vssio
port 624 nsew
flabel metal5 705730 397828 706000 399878 0 FreeSans 1600 90 0 0 vssio
port 624 nsew
flabel metal5 705730 400198 706000 402248 0 FreeSans 1600 90 0 0 vssio
port 624 nsew
flabel metal5 705730 402828 706000 404728 0 FreeSans 1600 90 0 0 vssio
port 624 nsew
flabel metal5 705730 433272 706000 435172 0 FreeSans 1600 90 0 0 vssd
port 625 nsew
flabel metal5 705730 435752 706000 437802 0 FreeSans 1600 90 0 0 vssd
port 625 nsew
flabel metal5 705730 438122 706000 440172 0 FreeSans 1600 90 0 0 vssd
port 625 nsew
flabel metal5 705730 440828 706000 442878 0 FreeSans 1600 90 0 0 vssd
port 625 nsew
flabel metal5 705730 443198 706000 445248 0 FreeSans 1600 90 0 0 vssd
port 625 nsew
flabel metal5 705730 445828 706000 447728 0 FreeSans 1600 90 0 0 vssd
port 625 nsew
flabel metal5 705730 476272 706000 478172 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 705730 478752 706000 480802 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 705730 481122 706000 483172 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 705730 483828 706000 485878 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 705730 486198 706000 488248 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 705730 488828 706000 490728 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 705726 777248 706004 779196 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 705730 779752 706000 781802 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 705728 782110 706002 784184 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 705730 784828 706000 786878 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 705728 787186 706002 789260 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 705730 789828 706000 791728 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 705728 863260 706002 865184 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 705730 865752 706000 867802 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 705728 868110 706002 870184 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 705730 870828 706000 872878 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 705728 873186 706002 875260 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 705730 875828 706000 877728 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 70000 85272 70270 87172 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 69998 87740 70272 89814 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 70000 90122 70270 92172 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 70000 92828 70270 94878 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 69998 95186 70272 97260 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 70000 97828 70270 99728 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 70000 126272 70270 128172 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 69998 128740 70272 130814 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 131122 70270 133172 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 133828 70270 135878 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 69998 136186 70272 138260 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 138828 70270 140728 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 413272 70270 415172 0 FreeSans 1600 90 0 0 vssd
port 625 nsew
flabel metal5 69998 415740 70272 417814 0 FreeSans 1600 90 0 0 vssd
port 625 nsew
flabel metal5 70000 418122 70270 420172 0 FreeSans 1600 90 0 0 vssd
port 625 nsew
flabel metal5 70000 420828 70270 422878 0 FreeSans 1600 90 0 0 vssd
port 625 nsew
flabel metal5 69998 423186 70272 425260 0 FreeSans 1600 90 0 0 vssd
port 625 nsew
flabel metal5 70000 425828 70270 427728 0 FreeSans 1600 90 0 0 vssd
port 625 nsew
flabel metal5 70000 454272 70270 456172 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 456752 70270 458802 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 459122 70270 461172 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 461828 70270 463878 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 464198 70270 466248 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 466828 70270 468728 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 782273 70270 784173 0 FreeSans 1600 90 0 0 vssio
port 624 nsew
flabel metal5 70000 784753 70270 786803 0 FreeSans 1600 90 0 0 vssio
port 624 nsew
flabel metal5 70000 787123 70270 789173 0 FreeSans 1600 90 0 0 vssio
port 624 nsew
flabel metal5 70000 789829 70270 791879 0 FreeSans 1600 90 0 0 vssio
port 624 nsew
flabel metal5 70000 792199 70270 794249 0 FreeSans 1600 90 0 0 vssio
port 624 nsew
flabel metal5 70000 794829 70270 796729 0 FreeSans 1600 90 0 0 vssio
port 624 nsew
flabel metal5 70000 823272 70270 825172 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 825752 70270 827802 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 828122 70270 830172 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 830828 70270 832878 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 833198 70270 835248 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 835828 70270 837728 0 FreeSans 1600 90 0 0 vddio
port 626 nsew
flabel metal5 70000 864272 70270 866172 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 70000 866752 70270 868802 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 70000 869122 70270 871172 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 70000 871828 70270 873878 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 70000 874198 70270 876248 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal5 70000 876828 70270 878728 0 FreeSans 1600 90 0 0 vccd
port 627 nsew
flabel metal2 162066 69900 162142 70200 0 FreeSans 480 90 0 0 resetb_pulldown
port 586 nsew
flabel metal3 705729 104558 706029 104634 0 FreeSans 480 0 0 0 gpio_loopback_one[0]
port 497 nsew
flabel metal3 705729 104746 706029 104822 0 FreeSans 480 0 0 0 gpio_loopback_zero[0]
port 496 nsew
flabel metal3 705729 147558 706029 147634 0 FreeSans 480 0 0 0 gpio_loopback_one[1]
port 499 nsew
flabel metal3 705729 147746 706029 147822 0 FreeSans 480 0 0 0 gpio_loopback_zero[1]
port 498 nsew
flabel metal3 705729 190558 706029 190634 0 FreeSans 480 0 0 0 gpio_loopback_one[2]
port 501 nsew
flabel metal3 705729 190746 706029 190822 0 FreeSans 480 0 0 0 gpio_loopback_zero[2]
port 500 nsew
flabel metal3 705729 233746 706029 233822 0 FreeSans 480 0 0 0 gpio_loopback_zero[3]
port 503 nsew
flabel metal3 705729 233558 706029 233634 0 FreeSans 480 0 0 0 gpio_loopback_one[3]
port 502 nsew
flabel metal3 705729 319746 706029 319822 0 FreeSans 480 0 0 0 gpio_loopback_zero[5]
port 507 nsew
flabel metal3 705729 319558 706029 319634 0 FreeSans 480 0 0 0 gpio_loopback_one[5]
port 506 nsew
flabel metal3 705729 534746 706029 534822 0 FreeSans 480 0 0 0 gpio_loopback_zero[7]
port 511 nsew
flabel metal3 705729 534558 706029 534634 0 FreeSans 480 0 0 0 gpio_loopback_one[7]
port 510 nsew
flabel metal3 705729 620746 706029 620822 0 FreeSans 480 0 0 0 gpio_loopback_zero[9]
port 515 nsew
flabel metal3 705729 620558 706029 620634 0 FreeSans 480 0 0 0 gpio_loopback_one[9]
port 514 nsew
flabel metal3 705729 706746 706029 706822 0 FreeSans 480 0 0 0 gpio_loopback_zero[11]
port 519 nsew
flabel metal3 705729 706558 706029 706634 0 FreeSans 480 0 0 0 gpio_loopback_one[11]
port 518 nsew
flabel metal3 705729 749558 706029 749634 0 FreeSans 480 0 0 0 gpio_loopback_one[12]
port 521 nsew
flabel metal3 705729 749746 706029 749822 0 FreeSans 480 0 0 0 gpio_loopback_zero[12]
port 520 nsew
flabel metal3 705729 921558 706029 921634 0 FreeSans 480 0 0 0 gpio_loopback_one[14]
port 525 nsew
flabel metal3 705729 921746 706029 921822 0 FreeSans 480 0 0 0 gpio_loopback_zero[14]
port 524 nsew
flabel metal3 705729 276558 706029 276634 0 FreeSans 480 0 0 0 gpio_loopback_one[4]
port 505 nsew
flabel metal3 705729 276746 706029 276822 0 FreeSans 480 0 0 0 gpio_loopback_zero[4]
port 504 nsew
flabel metal3 705729 362558 706029 362634 0 FreeSans 480 0 0 0 gpio_loopback_one[6]
port 509 nsew
flabel metal3 705729 362746 706029 362822 0 FreeSans 480 0 0 0 gpio_loopback_zero[6]
port 508 nsew
flabel metal3 705729 577746 706029 577822 0 FreeSans 480 0 0 0 gpio_loopback_zero[8]
port 512 nsew
flabel metal3 705729 577558 706029 577634 0 FreeSans 480 0 0 0 gpio_loopback_one[8]
port 513 nsew
flabel metal3 705729 663746 706029 663822 0 FreeSans 480 0 0 0 gpio_loopback_zero[10]
port 516 nsew
flabel metal3 705729 663558 706029 663634 0 FreeSans 480 0 0 0 gpio_loopback_one[10]
port 517 nsew
flabel metal3 705729 835746 706029 835822 0 FreeSans 480 0 0 0 gpio_loopback_zero[13]
port 523 nsew
flabel metal3 705729 835558 706029 835634 0 FreeSans 480 0 0 0 gpio_loopback_one[13]
port 522 nsew
flabel metal2 653178 943800 653254 944100 0 FreeSans 480 90 0 0 gpio_loopback_zero[15]
port 527 nsew
flabel metal2 653366 943800 653442 944100 0 FreeSans 480 90 0 0 gpio_loopback_one[15]
port 526 nsew
flabel metal2 543178 943800 543254 944100 0 FreeSans 480 90 0 0 gpio_loopback_zero[16]
port 528 nsew
flabel metal2 543366 943800 543442 944100 0 FreeSans 480 90 0 0 gpio_loopback_one[16]
port 529 nsew
flabel metal2 433178 943800 433254 944100 0 FreeSans 480 90 0 0 gpio_loopback_zero[18]
port 532 nsew
flabel metal2 433366 943800 433442 944100 0 FreeSans 480 90 0 0 gpio_loopback_one[18]
port 533 nsew
flabel metal2 268178 943800 268254 944100 0 FreeSans 480 90 0 0 gpio_loopback_zero[20]
port 536 nsew
flabel metal2 268366 943800 268442 944100 0 FreeSans 480 90 0 0 gpio_loopback_one[20]
port 537 nsew
flabel metal2 158178 943800 158254 944100 0 FreeSans 480 90 0 0 gpio_loopback_zero[22]
port 540 nsew
flabel metal2 158366 943800 158442 944100 0 FreeSans 480 90 0 0 gpio_loopback_one[22]
port 541 nsew
flabel metal3 69971 904178 70271 904254 0 FreeSans 480 0 0 0 gpio_loopback_zero[24]
port 544 nsew
flabel metal3 69971 740366 70271 740442 0 FreeSans 480 0 0 0 gpio_loopback_one[25]
port 546 nsew
flabel metal3 69971 740178 70271 740254 0 FreeSans 480 0 0 0 gpio_loopback_zero[25]
port 547 nsew
flabel metal3 69971 658178 70271 658254 0 FreeSans 480 0 0 0 gpio_loopback_zero[27]
port 551 nsew
flabel metal3 69971 658366 70271 658442 0 FreeSans 480 0 0 0 gpio_loopback_one[27]
port 550 nsew
flabel metal3 69971 576178 70271 576254 0 FreeSans 480 0 0 0 gpio_loopback_zero[29]
port 555 nsew
flabel metal3 69971 576366 70271 576442 0 FreeSans 480 0 0 0 gpio_loopback_one[29]
port 554 nsew
flabel metal3 69971 494178 70271 494254 0 FreeSans 480 0 0 0 gpio_loopback_zero[31]
port 559 nsew
flabel metal3 69971 494366 70271 494442 0 FreeSans 480 0 0 0 gpio_loopback_one[31]
port 558 nsew
flabel metal3 69971 371366 70271 371442 0 FreeSans 480 0 0 0 gpio_loopback_one[32]
port 561 nsew
flabel metal3 69971 330178 70271 330254 0 FreeSans 480 0 0 0 gpio_loopback_zero[33]
port 563 nsew
flabel metal3 69971 330366 70271 330442 0 FreeSans 480 0 0 0 gpio_loopback_one[33]
port 562 nsew
flabel metal3 69971 289366 70271 289442 0 FreeSans 480 0 0 0 gpio_loopback_one[34]
port 565 nsew
flabel metal3 69972 248178 70271 248254 0 FreeSans 480 0 0 0 gpio_loopback_zero[35]
port 567 nsew
flabel metal3 69972 248366 70271 248442 0 FreeSans 480 0 0 0 gpio_loopback_one[35]
port 566 nsew
flabel metal3 69971 207366 70271 207442 0 FreeSans 480 0 0 0 gpio_loopback_one[36]
port 569 nsew
flabel metal3 69971 166178 70271 166254 0 FreeSans 480 0 0 0 gpio_loopback_zero[37]
port 571 nsew
flabel metal3 69971 166366 70271 166442 0 FreeSans 480 0 0 0 gpio_loopback_one[37]
port 570 nsew
flabel metal2 340746 69900 340822 70200 0 FreeSans 480 90 0 0 gpio_loopback_zero[39]
port 576 nsew
flabel metal2 340558 69900 340634 70200 0 FreeSans 480 90 0 0 gpio_loopback_one[39]
port 574 nsew
flabel metal2 450746 69900 450822 70200 0 FreeSans 480 90 0 0 gpio_loopback_zero[41]
port 580 nsew
flabel metal2 450558 69900 450634 70200 0 FreeSans 480 90 0 0 gpio_loopback_one[41]
port 579 nsew
flabel metal2 560746 69900 560822 70200 0 FreeSans 480 90 0 0 gpio_loopback_zero[43]
port 584 nsew
flabel metal2 560558 69900 560634 70200 0 FreeSans 480 90 0 0 gpio_loopback_one[43]
port 583 nsew
flabel metal2 161194 69900 161270 70200 0 FreeSans 480 90 0 0 resetb_pullup
port 585 nsew
<< properties >>
string FIXED_BBOX 70017 70017 705983 943983
<< end >>
